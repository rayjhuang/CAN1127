
module chiptop_1127a0 ( CSP, CSN, VFB, COM, LG, SW, HG, BST, GATE, VDRV, DP, 
        DN, CC1, CC2, TST, GPIO_TS, SCL, SDA, GPIO1, GPIO2, GPIO3, GPIO4, 
        GPIO5 );
  input TST;
  inout CSP,  CSN,  VFB,  COM,  LG,  SW,  HG,  BST,  GATE,  VDRV,  DP,  DN, 
     CC1,  CC2,  GPIO_TS,  SCL,  SDA,  GPIO1,  GPIO2,  GPIO3,  GPIO4,  GPIO5;
  wire   SRAM_WEB, SRAM_CEB, SRAM_OEB, RD_ENB, STB_RP, DRP_OSC, IMP_OSC, TX_EN,
         TX_DAT, RX_DAT, RX_SQL, DAC1_EN, AD_RST, AD_HOLD, COMP_O, CCI2C_EN,
         RSTB, SLEEP, OSC_LOW, OSC_STOP, PWRDN, VPP_0V, VPP_SEL, LDO3P9V,
         OSC_O, RD_DET, OCP_SEL, CC1_DOB, CC2_DOB, CC1_DI, CC2_DI, DP_COMP,
         DN_COMP, DN_FAULT, PWREN_HOLD, LFOSC_ENB, VPP_OTP, IO_RSTB5, V1P1,
         ANAP_TS, TS_ANA_R, ANAP_GP1, GP1_ANA_R, ANAP_GP2, GP2_ANA_R, ANAP_GP3,
         GP3_ANA_R, ANAP_GP4, GP4_ANA_R, ANAP_GP5, GP5_ANA_R, DI_TST, DI_TS,
         SRAM_CLK, PMEM_RE, PMEM_PGM, PMEM_CSB, do_ccctl_0_, do_srcctl_0,
         tm_atpg, SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2,
         SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4,
         SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6,
         SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8,
         SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10,
         SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12,
         SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14,
         SYNOPSYS_UNCONNECTED_15, SYNOPSYS_UNCONNECTED_16,
         SYNOPSYS_UNCONNECTED_17, SYNOPSYS_UNCONNECTED_18,
         SYNOPSYS_UNCONNECTED_19, SYNOPSYS_UNCONNECTED_20,
         SYNOPSYS_UNCONNECTED_21, SYNOPSYS_UNCONNECTED_22,
         SYNOPSYS_UNCONNECTED_23, SYNOPSYS_UNCONNECTED_24,
         SYNOPSYS_UNCONNECTED_25;
  wire   [10:0] SRAM_A;
  wire   [7:0] SRAM_D;
  wire   [7:0] ANAOPT;
  wire   [1:0] FSW;
  wire   [1:0] RP_EN;
  wire   [1:0] VCONN_EN;
  wire   [17:0] SAMPL_SEL;
  wire   [7:0] DUMMY_IN;
  wire   [55:0] REGTRM;
  wire   [7:0] PWR_I;
  wire   [1:0] OVP_SEL;
  wire   [5:0] DAC3_V;
  wire   [10:0] DAC0;
  wire   [3:0] ANA_TM;
  wire   [9:0] DAC1;
  wire   [1:0] RP_SEL;
  wire   [1:0] IE_GPIO;
  wire   [6:0] DI_GPIO;
  wire   [6:0] OE_GPIO;
  wire   [6:0] DO_GPIO;
  wire   [6:0] PU_GPIO;
  wire   [6:0] PD_GPIO;
  wire   [3:0] DO_TS;
  wire   [1:0] PMEM_CLK;
  wire   [7:0] PMEM_Q1;
  wire   [7:0] PMEM_Q0;
  wire   [1:0] PMEM_SAP;
  wire   [1:0] PMEM_TWLB;
  wire   [15:0] PMEM_A;
  wire   [6:0] bck_regx0;
  wire   [7:2] do_xana1;
  wire   [7:0] do_xana0;
  wire   [3:0] do_regx_xtm;
  wire   [5:2] do_cvctl;
  wire   [3:0] do_vooc;
  wire   [5:0] do_dpdm;
  wire   [5:4] do_srcctl;
  wire   [7:0] do_cctrx;
  wire   [3:0] di_xanav;
  wire   [5:0] srci;
  tri   VFB;
  tri   COM;
  tri   LG;
  tri   SW;
  tri   HG;
  tri   BST;
  tri   GATE;
  tri   VDRV;
  tri   DP;
  tri   DN;
  tri   CC1;
  tri   CC2;
  tri   TST;
  tri   GPIO_TS;
  tri   SCL;
  tri   SDA;
  tri   GPIO1;
  tri   GPIO2;
  tri   GPIO3;
  tri   GPIO4;
  tri   GPIO5;
  tri   [7:0] xdat_o;

  anatop_1127a0 U0_ANALOG_TOP ( .CC1(CC1), .CC2(CC2), .DP(DP), .DN(DN), .VFB(
        VFB), .CSP(), .CSN(), .COM(COM), .LG(LG), .SW(SW), .HG(HG), .BST(BST), 
        .GATE(GATE), .VDRV(VDRV), .BST_SET(bck_regx0[0]), .DCM_SEL(
        bck_regx0[1]), .HGOFF(bck_regx0[2]), .HGLGOFF(bck_regx0[3]), .HGON(
        bck_regx0[4]), .LGON(bck_regx0[5]), .ENDRV(bck_regx0[6]), .FSW(FSW), 
        .EN_OSC(bck_regx0[2]), .MAXDS(bck_regx0[3]), .EN_GM(bck_regx0[4]), 
        .EN_ODLDO(bck_regx0[5]), .EN_IBUK(bck_regx0[6]), .RP_SEL(RP_SEL), 
        .RP1_EN(RP_EN[0]), .RP2_EN(RP_EN[1]), .VCONN1_EN(VCONN_EN[0]), 
        .VCONN2_EN(VCONN_EN[1]), .SGP({do_cctrx[0], do_regx_xtm}), .S20U(
        do_cctrx[1]), .S100U(do_cctrx[2]), .TX_EN(TX_EN), .TX_DAT(TX_DAT), 
        .CC_SEL(do_ccctl_0_), .TRA(do_cctrx[4]), .TFA(do_cctrx[5]), .LSR(
        do_cctrx[6]), .RX_DAT(RX_DAT), .RX_SQL(RX_SQL), .SEL_RX_TH(do_cctrx[7]), .DAC1_EN(DAC1_EN), .DPDN_SHORT(do_dpdm[0]), .DP_2V7_EN(do_dpdm[4]), 
        .DN_2V7_EN(do_dpdm[3]), .DP_0P6V_EN(do_xana1[3]), .DN_0P6V_EN(
        do_xana1[2]), .DP_DWN_EN(do_dpdm[2]), .DN_DWN_EN(do_dpdm[1]), .PWR_I(
        PWR_I), .DAC3(DAC3_V), .DAC1(DAC1), .CV2(do_xana0[0]), .LFOSC_ENB(
        LFOSC_ENB), .VO_DISCHG(do_srcctl[4]), .DISCHG_SEL(do_srcctl[5]), 
        .CMP_SEL_VO10(SAMPL_SEL[0]), .CMP_SEL_VO20(SAMPL_SEL[10]), 
        .CMP_SEL_GP1(SAMPL_SEL[17]), .CMP_SEL_GP2(SAMPL_SEL[16]), 
        .CMP_SEL_GP3(SAMPL_SEL[15]), .CMP_SEL_GP4(SAMPL_SEL[14]), 
        .CMP_SEL_GP5(SAMPL_SEL[13]), .CMP_SEL_VIN20(SAMPL_SEL[1]), 
        .CMP_SEL_TS(SAMPL_SEL[3]), .CMP_SEL_IS(SAMPL_SEL[2]), .CMP_SEL_CC2(
        SAMPL_SEL[7]), .CMP_SEL_CC1(SAMPL_SEL[6]), .CMP_SEL_CC2_4(
        SAMPL_SEL[12]), .CMP_SEL_CC1_4(SAMPL_SEL[11]), .CMP_SEL_DP(
        SAMPL_SEL[4]), .CMP_SEL_DP_3(SAMPL_SEL[8]), .CMP_SEL_DN(SAMPL_SEL[5]), 
        .CMP_SEL_DN_3(SAMPL_SEL[9]), .OCP_EN(do_cvctl[2]), .CS_EN(do_cctrx[3]), 
        .COMP_O(COMP_O), .CCI2C_EN(CCI2C_EN), .UVP_SEL(do_xana0[7]), .TM(
        ANA_TM), .V5OCP(srci[4]), .RSTB(RSTB), .DAC0(DAC0), .SLEEP(SLEEP), 
        .OSC_LOW(OSC_LOW), .OSC_STOP(OSC_STOP), .PWRDN(PWRDN), .VPP_ZERO(
        VPP_0V), .OSC_O(OSC_O), .RD_DET(RD_DET), .IMP_OSC(IMP_OSC), .DRP_OSC(
        DRP_OSC), .STB_RP(STB_RP), .RD_ENB(RD_ENB), .PWREN(do_srcctl_0), .OCP(
        srci[1]), .SCP(srci[3]), .UVP(srci[0]), .LDO3P9V(LDO3P9V), .VPP_SEL(
        VPP_SEL), .CC1_DOB(CC1_DOB), .CC2_DOB(CC2_DOB), .CC1_DI(CC1_DI), 
        .CC2_DI(CC2_DI), .ANTI_INRUSH(do_cvctl[5]), .OTPI(srci[5]), .OVP_SEL(
        OVP_SEL), .OVP(srci[2]), .DN_COMP(DN_COMP), .DP_COMP(DP_COMP), 
        .DPDN_VTH(do_xana0[5]), .DPDEN(do_vooc[3]), .DPDO(do_vooc[2]), .DPIE(
        do_dpdm[5]), .DNDEN(do_vooc[1]), .DNDO(do_vooc[0]), .DNIE(do_dpdm[5]), 
        .DUMMY_IN(DUMMY_IN), .CP_CLKX2(ANAOPT[7]), .SEL_CONST_OVP(ANAOPT[6]), 
        .LP_EN(ANAOPT[5]), .DNCHK_EN(ANAOPT[3]), .IRP_EN(ANAOPT[2]), .CCBFEN(
        ANAOPT[0]), .REGTRM(REGTRM), .AD_RST(AD_RST), .AD_HOLD(AD_HOLD), 
        .DN_FAULT(DN_FAULT), .SEL_CCGAIN(do_xana0[3]), .VFB_SW(do_xana0[1]), 
        .CPV_SEL(do_xana1[6]), .CLAMPV_EN(do_xana1[5]), .HVNG_CPEN(do_xana1[7]), .PWREN_HOLD(PWREN_HOLD), .OCP_SEL(OCP_SEL), .OCP_80M(di_xanav[1]), 
        .OCP_160M(di_xanav[0]), .OPTO1(di_xanav[2]), .OPTO2(di_xanav[3]), 
        .VPP_OTP(VPP_OTP), .VDD_OTP(), .RSTB_5(IO_RSTB5), .V1P1(V1P1), 
        .TS_ANA_R(TS_ANA_R), .GP5_ANA_R(GP5_ANA_R), .GP4_ANA_R(GP4_ANA_R), 
        .GP3_ANA_R(GP3_ANA_R), .GP2_ANA_R(GP2_ANA_R), .GP1_ANA_R(GP1_ANA_R), 
        .TS_ANA_P(ANAP_TS), .GP5_ANA_P(ANAP_GP5), .GP4_ANA_P(ANAP_GP4), 
        .GP3_ANA_P(ANAP_GP3), .GP2_ANA_P(ANAP_GP2), .GP1_ANA_P(ANAP_GP1) );
  IODMURUDA_A0 PAD_SCL ( .DO(DO_GPIO[0]), .IE(IE_GPIO[1]), .OE(OE_GPIO[0]), 
        .PD(PD_GPIO[0]), .PU(PU_GPIO[0]), .RSTB_5(IO_RSTB5), .VB(V1P1), .PAD(
        SCL), .ANA_R(), .DI(DI_GPIO[0]) );
  IODMURUDA_A0 PAD_SDA ( .DO(DO_GPIO[1]), .IE(IE_GPIO[1]), .OE(OE_GPIO[1]), 
        .PD(PD_GPIO[1]), .PU(PU_GPIO[1]), .RSTB_5(IO_RSTB5), .VB(V1P1), .PAD(
        SDA), .ANA_R(), .DI(DI_GPIO[1]) );
  IOBMURUDA_A0 PAD_TST ( .DO(1'b0), .IE(1'b1), .OE(1'b0), .PD(1'b1), .PU(1'b0), 
        .RSTB_5(IO_RSTB5), .VB(V1P1), .PAD(TST), .ANA_R(), .DI(DI_TST) );
  IOBMURUDA_A1 PAD_GPIO1 ( .ANA_P(ANAP_GP1), .DO(DO_GPIO[2]), .IE(IE_GPIO[0]), 
        .OE(OE_GPIO[2]), .PD(PD_GPIO[2]), .PU(PU_GPIO[2]), .RSTB_5(IO_RSTB5), 
        .VB(V1P1), .PAD(GPIO1), .ANA_R(GP1_ANA_R), .DI(DI_GPIO[2]) );
  IOBMURUDA_A1 PAD_GPIO2 ( .ANA_P(ANAP_GP2), .DO(DO_GPIO[3]), .IE(IE_GPIO[0]), 
        .OE(OE_GPIO[3]), .PD(PD_GPIO[3]), .PU(PU_GPIO[3]), .RSTB_5(IO_RSTB5), 
        .VB(V1P1), .PAD(GPIO2), .ANA_R(GP2_ANA_R), .DI(DI_GPIO[3]) );
  IOBMURUDA_A1 PAD_GPIO3 ( .ANA_P(ANAP_GP3), .DO(DO_GPIO[4]), .IE(IE_GPIO[0]), 
        .OE(OE_GPIO[4]), .PD(PD_GPIO[4]), .PU(PU_GPIO[4]), .RSTB_5(IO_RSTB5), 
        .VB(V1P1), .PAD(GPIO3), .ANA_R(GP3_ANA_R), .DI(DI_GPIO[4]) );
  IOBMURUDA_A1 PAD_GPIO4 ( .ANA_P(ANAP_GP4), .DO(DO_GPIO[5]), .IE(IE_GPIO[0]), 
        .OE(OE_GPIO[5]), .PD(PD_GPIO[5]), .PU(PU_GPIO[5]), .RSTB_5(IO_RSTB5), 
        .VB(V1P1), .PAD(GPIO4), .ANA_R(GP4_ANA_R), .DI(DI_GPIO[5]) );
  IOBMURUDA_A1 PAD_GPIO5 ( .ANA_P(ANAP_GP5), .DO(DO_GPIO[6]), .IE(IE_GPIO[0]), 
        .OE(OE_GPIO[6]), .PD(PD_GPIO[6]), .PU(PU_GPIO[6]), .RSTB_5(IO_RSTB5), 
        .VB(V1P1), .PAD(GPIO5), .ANA_R(GP5_ANA_R), .DI(DI_GPIO[6]) );
  IOBMURUDA_A1 PAD_GPIO_TS ( .ANA_P(ANAP_TS), .DO(DO_TS[3]), .IE(IE_GPIO[0]), 
        .OE(DO_TS[2]), .PD(DO_TS[0]), .PU(DO_TS[1]), .RSTB_5(IO_RSTB5), .VB(
        V1P1), .PAD(GPIO_TS), .ANA_R(TS_ANA_R), .DI(DI_TS) );
  MSL18B_1536X8_RW10TM4_16 U0_SRAM ( .A(SRAM_A), .DI(SRAM_D), .DO(xdat_o), 
        .CK(SRAM_CLK), .WEB(SRAM_WEB), .CSB(SRAM_CEB), .OEB(SRAM_OEB) );
  ATO0008KX8MX180LBX4DA U0_CODE_0_ ( .A(PMEM_A), .TWLB(PMEM_TWLB), .Q(PMEM_Q0), 
        .SAP(PMEM_SAP), .CSB(PMEM_CSB), .CLK(PMEM_CLK[0]), .PGM(PMEM_PGM), 
        .RE(PMEM_RE), .VDDP(VPP_OTP), .VDD(), .VSS() );
  ATO0008KX8MX180LBX4DA U0_CODE_1_ ( .A(PMEM_A), .TWLB(PMEM_TWLB), .Q(PMEM_Q1), 
        .SAP(PMEM_SAP), .CSB(PMEM_CSB), .CLK(PMEM_CLK[1]), .PGM(PMEM_PGM), 
        .RE(PMEM_RE), .VDDP(VPP_OTP), .VDD(), .VSS() );
  core_a0 U0_CORE ( .SRCI(srci), .XANAV({1'b0, di_xanav}), .BCK_REGX({
        SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3, 
        SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6, 
        FSW, SYNOPSYS_UNCONNECTED_7, bck_regx0}), .ANA_REGX({do_xana1[7:5], 
        SYNOPSYS_UNCONNECTED_8, do_xana1[3:2], SYNOPSYS_UNCONNECTED_9, 
        SYNOPSYS_UNCONNECTED_10, do_xana0[7], SYNOPSYS_UNCONNECTED_11, 
        do_xana0[5], SYNOPSYS_UNCONNECTED_12, do_xana0[3], 
        SYNOPSYS_UNCONNECTED_13, do_xana0[1:0]}), .LFOSC_ENB(LFOSC_ENB), 
        .STB_RP(STB_RP), .RD_ENB(RD_ENB), .OCP_SEL(OCP_SEL), .PWREN_HOLD(
        PWREN_HOLD), .CC1_DI(CC1_DI), .CC2_DI(CC2_DI), .DRP_OSC(DRP_OSC), 
        .IMP_OSC(IMP_OSC), .CC1_DOB(CC1_DOB), .CC2_DOB(CC2_DOB), .DAC1_EN(
        DAC1_EN), .SH_RST(AD_RST), .SH_HOLD(AD_HOLD), .LDO3P9V(LDO3P9V), .XTM(
        do_regx_xtm), .DO_CVCTL({OVP_SEL, do_cvctl[5], SYNOPSYS_UNCONNECTED_14, 
        SYNOPSYS_UNCONNECTED_15, do_cvctl[2], SYNOPSYS_UNCONNECTED_16, 
        SYNOPSYS_UNCONNECTED_17}), .DO_CCTRX(do_cctrx), .DO_SRCCTL({
        SYNOPSYS_UNCONNECTED_18, SYNOPSYS_UNCONNECTED_19, do_srcctl, VCONN_EN, 
        SYNOPSYS_UNCONNECTED_20, do_srcctl_0}), .DO_CCCTL({RP_EN, RP_SEL, 
        SYNOPSYS_UNCONNECTED_21, SYNOPSYS_UNCONNECTED_22, 
        SYNOPSYS_UNCONNECTED_23, do_ccctl_0_}), .DO_DAC0(DAC0), .DO_DPDN(
        do_dpdm), .DO_VOOC(do_vooc), .DO_PWR_I(PWR_I), .PMEM_A(PMEM_A), 
        .PMEM_Q0(PMEM_Q0), .PMEM_Q1(PMEM_Q1), .PMEM_TWLB(PMEM_TWLB), 
        .PMEM_SAP(PMEM_SAP), .PMEM_CLK(PMEM_CLK), .PMEM_CSB(PMEM_CSB), 
        .PMEM_RE(PMEM_RE), .PMEM_PGM(PMEM_PGM), .VPP_SEL(VPP_SEL), .VPP_0V(
        VPP_0V), .SRAM_WEB(SRAM_WEB), .SRAM_CEB(SRAM_CEB), .SRAM_OEB(SRAM_OEB), 
        .SRAM_CLK(SRAM_CLK), .SRAM_A(SRAM_A), .SRAM_D(SRAM_D), .SRAM_RDAT(
        xdat_o), .RX_DAT(RX_DAT), .RX_SQL(RX_SQL), .RD_DET(RD_DET), .STB_OVP(
        1'b0), .TX_DAT(TX_DAT), .TX_EN(TX_EN), .OSC_STOP(OSC_STOP), .OSC_LOW(
        OSC_LOW), .SLEEP(SLEEP), .PWRDN(PWRDN), .OCDRV_ENZ(), .DAC1_V(DAC1), 
        .SAMPL_SEL(SAMPL_SEL), .DAC1_COMP(COMP_O), .CCI2C_EN(CCI2C_EN), 
        .ANA_TM(ANA_TM), .DM_FAULT(DN_FAULT), .DM_COMP(DN_COMP), .DP_COMP(
        DP_COMP), .DI_GPIO(DI_GPIO), .DO_GPIO(DO_GPIO), .OE_GPIO(OE_GPIO), 
        .GPIO_PU(PU_GPIO), .GPIO_PD(PD_GPIO), .GPIO_IE(IE_GPIO), .DO_TS(DO_TS), 
        .DI_TS(DI_TS), .REGTRM(REGTRM), .ANAOPT({ANAOPT[7:5], 
        SYNOPSYS_UNCONNECTED_24, ANAOPT[3:2], SYNOPSYS_UNCONNECTED_25, 
        ANAOPT[0]}), .DUMMY_IN(DUMMY_IN), .DAC3_V(DAC3_V), .i_clk(OSC_O), 
        .i_rstz(RSTB), .atpg_en(tm_atpg), .di_tst(DI_TST), .tm_atpg(tm_atpg)
         );
endmodule


module core_a0 ( SRCI, XANAV, BCK_REGX, ANA_REGX, LFOSC_ENB, STB_RP, RD_ENB, 
        OCP_SEL, PWREN_HOLD, CC1_DI, CC2_DI, DRP_OSC, IMP_OSC, CC1_DOB, 
        CC2_DOB, DAC1_EN, SH_RST, SH_HOLD, LDO3P9V, XTM, DO_CVCTL, DO_CCTRX, 
        DO_SRCCTL, DO_CCCTL, DO_DAC0, DO_DPDN, DO_VOOC, DO_PWR_I, PMEM_A, 
        PMEM_Q0, PMEM_Q1, PMEM_TWLB, PMEM_SAP, PMEM_CLK, PMEM_CSB, PMEM_RE, 
        PMEM_PGM, VPP_SEL, VPP_0V, SRAM_WEB, SRAM_CEB, SRAM_OEB, SRAM_CLK, 
        SRAM_A, SRAM_D, SRAM_RDAT, RX_DAT, RX_SQL, RD_DET, STB_OVP, TX_DAT, 
        TX_EN, OSC_STOP, OSC_LOW, SLEEP, PWRDN, OCDRV_ENZ, DAC1_V, SAMPL_SEL, 
        DAC1_COMP, CCI2C_EN, ANA_TM, DM_FAULT, DM_COMP, DP_COMP, DI_GPIO, 
        DO_GPIO, OE_GPIO, GPIO_PU, GPIO_PD, GPIO_IE, DO_TS, DI_TS, REGTRM, 
        ANAOPT, DUMMY_IN, DAC3_V, i_clk, i_rstz, atpg_en, di_tst, tm_atpg );
  input [5:0] SRCI;
  input [4:0] XANAV;
  output [15:0] BCK_REGX;
  output [15:0] ANA_REGX;
  output [3:0] XTM;
  output [7:0] DO_CVCTL;
  output [7:0] DO_CCTRX;
  output [7:0] DO_SRCCTL;
  output [7:0] DO_CCCTL;
  output [10:0] DO_DAC0;
  output [5:0] DO_DPDN;
  output [3:0] DO_VOOC;
  output [7:0] DO_PWR_I;
  output [15:0] PMEM_A;
  input [7:0] PMEM_Q0;
  input [7:0] PMEM_Q1;
  output [1:0] PMEM_TWLB;
  output [1:0] PMEM_SAP;
  output [1:0] PMEM_CLK;
  output [10:0] SRAM_A;
  output [7:0] SRAM_D;
  input [7:0] SRAM_RDAT;
  output [9:0] DAC1_V;
  output [17:0] SAMPL_SEL;
  output [3:0] ANA_TM;
  input [6:0] DI_GPIO;
  output [6:0] DO_GPIO;
  output [6:0] OE_GPIO;
  output [6:0] GPIO_PU;
  output [6:0] GPIO_PD;
  output [1:0] GPIO_IE;
  output [3:0] DO_TS;
  output [55:0] REGTRM;
  output [7:0] ANAOPT;
  output [7:0] DUMMY_IN;
  output [5:0] DAC3_V;
  input CC1_DI, CC2_DI, DRP_OSC, IMP_OSC, RX_DAT, RX_SQL, RD_DET, STB_OVP,
         DAC1_COMP, DM_FAULT, DM_COMP, DP_COMP, DI_TS, i_clk, i_rstz, atpg_en,
         di_tst;
  output LFOSC_ENB, STB_RP, RD_ENB, OCP_SEL, PWREN_HOLD, CC1_DOB, CC2_DOB,
         DAC1_EN, SH_RST, SH_HOLD, LDO3P9V, PMEM_CSB, PMEM_RE, PMEM_PGM,
         VPP_SEL, VPP_0V, SRAM_WEB, SRAM_CEB, SRAM_OEB, SRAM_CLK, TX_DAT,
         TX_EN, OSC_STOP, OSC_LOW, SLEEP, PWRDN, OCDRV_ENZ, CCI2C_EN, tm_atpg;
  wire   N258, N259, N260, N261, N262, N263, N264, N265, N266, N267, N268,
         N269, n626, n627, n628, n629, n630, aswclk, detclk, tclk_sel, s_clk,
         aswkup, x_clk, t_di_gpio4, r_osc_gate, g_clk, xram_ce, iram_ce,
         sram_en, r_i2c_attr, esfrm_oe, esfrm_we, sfrack, ictlr_psrack,
         esfrm_rrdy, memwr, memrd, memrd_c, memack, o_cpurst, hit_xd, hit_xr,
         hit_ps, hit_ps_c, mcu_ram_r, mcu_ram_w, regx_re, iram_we, xram_we,
         regx_we, bist_en, bist_wr, srstz, prl_cany0w, prl_cany0r, mempsrd,
         r_bclk_sel, r_hold_mcu, t0_intr, fcp_intr, dpdm_urx, s0_rxdoe,
         mcuo_scl, mcuo_sda, mempsack, mempswr, mempsrd_c, sfr_w, sfr_r,
         ictlr_psack, ictlr_inc, set_hold, bkpt_hold, bkpt_ena, r_psrd, r_pswr,
         prl_cany0, prl_c0set, pmem_pgm, pmem_re, pmem_csb, we_twlb,
         r_otp_wpls, pwrdn_rst, r_otp_pwdn_en, ramacc, r_sleep, ps_pwrdn,
         r_pwrdn, r_ocdrv_enz, r_osc_stop, r_pwrv_upd, r_otpi_gate, r_fcpre,
         r_fortxdat, r_fortxrdy, r_fortxen, r_gpio_tm, pid_goidle, pid_gobusy,
         bus_idle, sse_idle, r_exist1st, r_ordrs4, r_fifopsh, r_fifopop,
         r_unlock, r_first, r_last, r_fiforst, r_set_cpmsgid, r_txendk,
         r_txshrt, r_auto_discard, r_dat_portrole, r_dat_datarole, r_pshords,
         r_discard, r_strtch, r_i2c_ninc, r_i2c_fwnak, r_i2c_fwack,
         hwi2c_stretch, i2c_ev_6_, i2c_ev_3, i2c_ev_2, prl_discard,
         prl_GCTxDone, pff_obsd, pff_empty, pff_full, ptx_ack, clk_1500k,
         clk_500k, clk_500, prstz, sse_rdrdy, upd_rdrdy, sse_prefetch,
         slvo_sda, slvo_re, slvo_early, dm_comp, dp_comp, di_cc, ptx_cc,
         ptx_oe, sh_rst, sh_hold, fcp_oe, fcp_do, sdischg_duty, clk_100k,
         r_imp_osc, r_vpp_en, r_vpp0v_en, di_ts, r_xana_23, r_xana_19,
         r_xana_18, divff_8, divff_5, clk_50k, do_opt_1, do_opt_0, N449, N450,
         o_dodat0_15_, o_dodat5_2_, N570, N571, N572, N573, N574, N579, N580,
         N581, N582, N583, N584, N585, N586, N595, N596, N597, N598, N599,
         N600, N601, N602, N603, N604, N605, N606, N607, N608, N609, N610,
         N629, N630, N631, N632, N633, N634, N635, N636, N637, N638, N639,
         N640, N641, N642, N643, N644, N1483, N1488, N1493, N1498, net8831,
         n29, n30, n31, n77, n122, n124, n136, n138, n140, n142, n145, n147,
         n154, n156, n157, n158, n159, n160, n161, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n212, n213, n214, n215,
         n216, n217, n218, n220, n221, n222, n223, n224, n225, n226, n227,
         n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238,
         n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249,
         n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
         n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271,
         n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
         n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, sll_223_2_A_0_, n1, n2, n3, n4, n5, n6,
         n7, n9, n10, n11, n13, n14, n15, n16, n17, n18, n19, n23, n24, n25,
         n26, n27, n28, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n123, n125, n126, n127, n128, n129, n130, n131, n133, n134, n135,
         n137, n139, n141, n143, n144, n146, n148, n149, n150, n151, n152,
         n153, n155, n162, n163, n164, n165, n166, n211, n219, n508, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2,
         SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4,
         SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6,
         SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8,
         SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10,
         SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12,
         SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14,
         SYNOPSYS_UNCONNECTED_15, SYNOPSYS_UNCONNECTED_16,
         SYNOPSYS_UNCONNECTED_17, SYNOPSYS_UNCONNECTED_18,
         SYNOPSYS_UNCONNECTED_19, SYNOPSYS_UNCONNECTED_20,
         SYNOPSYS_UNCONNECTED_21, SYNOPSYS_UNCONNECTED_22,
         SYNOPSYS_UNCONNECTED_23, SYNOPSYS_UNCONNECTED_24,
         SYNOPSYS_UNCONNECTED_25, SYNOPSYS_UNCONNECTED_26,
         SYNOPSYS_UNCONNECTED_27, SYNOPSYS_UNCONNECTED_28,
         SYNOPSYS_UNCONNECTED_29, SYNOPSYS_UNCONNECTED_30,
         SYNOPSYS_UNCONNECTED_31, SYNOPSYS_UNCONNECTED_32,
         SYNOPSYS_UNCONNECTED_33, SYNOPSYS_UNCONNECTED_34,
         SYNOPSYS_UNCONNECTED_35, SYNOPSYS_UNCONNECTED_36,
         SYNOPSYS_UNCONNECTED_37, SYNOPSYS_UNCONNECTED_38,
         SYNOPSYS_UNCONNECTED_39, SYNOPSYS_UNCONNECTED_40,
         SYNOPSYS_UNCONNECTED_41, SYNOPSYS_UNCONNECTED_42,
         SYNOPSYS_UNCONNECTED_43, SYNOPSYS_UNCONNECTED_44,
         SYNOPSYS_UNCONNECTED_45, SYNOPSYS_UNCONNECTED_46,
         SYNOPSYS_UNCONNECTED_47, SYNOPSYS_UNCONNECTED_48,
         SYNOPSYS_UNCONNECTED_49, SYNOPSYS_UNCONNECTED_50,
         SYNOPSYS_UNCONNECTED_51, SYNOPSYS_UNCONNECTED_52,
         SYNOPSYS_UNCONNECTED_53, SYNOPSYS_UNCONNECTED_54,
         SYNOPSYS_UNCONNECTED_55, SYNOPSYS_UNCONNECTED_56,
         SYNOPSYS_UNCONNECTED_57, SYNOPSYS_UNCONNECTED_58,
         SYNOPSYS_UNCONNECTED_59, SYNOPSYS_UNCONNECTED_60,
         SYNOPSYS_UNCONNECTED_61, SYNOPSYS_UNCONNECTED_62,
         SYNOPSYS_UNCONNECTED_63, SYNOPSYS_UNCONNECTED_64,
         SYNOPSYS_UNCONNECTED_65, SYNOPSYS_UNCONNECTED_66,
         SYNOPSYS_UNCONNECTED_67, SYNOPSYS_UNCONNECTED_68,
         SYNOPSYS_UNCONNECTED_69, SYNOPSYS_UNCONNECTED_70,
         SYNOPSYS_UNCONNECTED_71, SYNOPSYS_UNCONNECTED_72,
         SYNOPSYS_UNCONNECTED_73, SYNOPSYS_UNCONNECTED_74,
         SYNOPSYS_UNCONNECTED_75, SYNOPSYS_UNCONNECTED_76,
         SYNOPSYS_UNCONNECTED_77, SYNOPSYS_UNCONNECTED_78,
         SYNOPSYS_UNCONNECTED_79, SYNOPSYS_UNCONNECTED_80,
         SYNOPSYS_UNCONNECTED_81, SYNOPSYS_UNCONNECTED_82,
         SYNOPSYS_UNCONNECTED_83, SYNOPSYS_UNCONNECTED_84,
         SYNOPSYS_UNCONNECTED_85, SYNOPSYS_UNCONNECTED_86,
         SYNOPSYS_UNCONNECTED_87, SYNOPSYS_UNCONNECTED_88,
         SYNOPSYS_UNCONNECTED_89, SYNOPSYS_UNCONNECTED_90,
         SYNOPSYS_UNCONNECTED_91, SYNOPSYS_UNCONNECTED_92,
         SYNOPSYS_UNCONNECTED_93, SYNOPSYS_UNCONNECTED_94,
         SYNOPSYS_UNCONNECTED_95, SYNOPSYS_UNCONNECTED_96,
         SYNOPSYS_UNCONNECTED_97, SYNOPSYS_UNCONNECTED_98,
         SYNOPSYS_UNCONNECTED_99, SYNOPSYS_UNCONNECTED_100,
         SYNOPSYS_UNCONNECTED_101;
  wire   [9:0] aswclk_ps;
  wire   [9:0] detclk_ps;
  wire   [7:0] sse_wdat;
  wire   [7:0] prx_fifowdat;
  wire   [7:0] sse_adr;
  wire   [7:0] prl_cany0adr;
  wire   [7:0] esfrm_wdat;
  wire   [6:0] esfrm_adr;
  wire   [7:0] mcu_esfrrdat;
  wire   [7:0] delay_inst;
  wire   [7:0] esfrm_rdat;
  wire   [3:0] r_pg0_sel;
  wire   [15:0] memaddr;
  wire   [15:0] memaddr_c;
  wire   [7:0] memdatao;
  wire   [7:0] idat_adr;
  wire   [7:0] idat_wdat;
  wire   [10:0] iram_a;
  wire   [10:0] xram_a;
  wire   [7:0] iram_d;
  wire   [7:0] xram_d;
  wire   [1:0] sram_rdat;
  wire   [7:0] regx_rdat;
  wire   [10:0] bist_adr;
  wire   [7:0] bist_wdat;
  wire   [7:0] memdatai;
  wire   [7:0] ictlr_inst;
  wire   [15:0] mcu_pc;
  wire   [22:16] mcu_dbgpo;
  wire   [3:2] sfr_intr;
  wire   [7:0] exint;
  wire   [7:0] ff_p0;
  wire   [6:0] do_p0;
  wire   [7:0] sfr_rdat;
  wire   [7:0] sfr_wdat;
  wire   [6:0] sfr_adr;
  wire   [14:0] bkpt_pc;
  wire   [14:0] r_inst_ofs;
  wire   [1:0] pmem_clk;
  wire   [7:0] pmem_q0;
  wire   [7:0] pmem_q1;
  wire   [1:0] pmem_twlb;
  wire   [1:0] wd_twlb;
  wire   [1:0] r_sqlch;
  wire   [3:2] r_ccrx;
  wire   [1:0] r_rxdb_opt;
  wire   [7:4] r_pwrctl;
  wire   [5:0] di_pro;
  wire   [7:0] r_cvctl;
  wire   [7:0] r_srcctl;
  wire   [7:0] r_dpdmctl;
  wire   [11:0] r_fw_pwrv;
  wire   [5:0] r_cvcwr;
  wire   [15:0] r_cvofs;
  wire   [7:0] r_cctrx;
  wire   [7:0] r_ccctl;
  wire   [6:0] r_fcpwr;
  wire   [7:0] fcp_r_dat;
  wire   [7:0] fcp_r_sta;
  wire   [7:0] fcp_r_msk;
  wire   [7:0] fcp_r_ctl;
  wire   [7:0] fcp_r_crc;
  wire   [7:0] fcp_r_acc;
  wire   [7:0] fcp_r_tui;
  wire   [7:0] r_accctl;
  wire   [7:5] r_comp_opt;
  wire   [14:0] sfr_dacwr;
  wire   [17:0] r_dac_en;
  wire   [17:0] r_sar_en;
  wire   [7:0] r_isofs;
  wire   [7:0] r_adofs;
  wire   [7:0] dac_r_ctl;
  wire   [7:0] dac_r_cmpsta;
  wire   [17:0] dac_r_comp;
  wire   [143:0] dac_r_vs;
  wire   [5:0] x_daclsb;
  wire   [6:0] REVID;
  wire   [6:0] r_pu_gpio;
  wire   [6:0] r_pd_gpio;
  wire   [6:0] r_gpio_oe;
  wire   [1:0] r_gpio_ie;
  wire   [55:0] r_regtrm;
  wire   [3:0] r_ana_tm;
  wire   [7:0] i2c_ltbuf;
  wire   [7:0] i2c_lt_ofs;
  wire   [4:0] r_txnumk;
  wire   [1:0] r_auto_gdcrc;
  wire   [1:0] r_spec;
  wire   [1:0] r_dat_spec;
  wire   [6:0] r_txauto;
  wire   [6:0] r_rxords_ena;
  wire   [7:1] r_i2c_deva;
  wire   [2:0] prl_cpmsgid;
  wire   [1:0] pff_ack;
  wire   [7:0] pff_rdat;
  wire   [15:0] pff_rxpart;
  wire   [5:0] pff_ptr;
  wire   [6:0] prx_setsta;
  wire   [1:0] prx_rst;
  wire   [4:0] prx_rcvinf;
  wire   [5:0] prx_adpn;
  wire   [3:0] prx_fsm;
  wire   [2:0] ptx_fsm;
  wire   [3:0] prl_fsm;
  wire   [3:0] slvo_ev;
  wire   [1:0] r_i2cslv_route;
  wire   [5:4] r_i2crout;
  wire   [1:0] r_i2cmcu_route;
  wire   [18:17] upd_dbgpo;
  wire   [7:0] r_dacwdat;
  wire   [17:8] wr_dacv;
  wire   [10:7] r_dacwr;
  wire   [17:0] dacmux_sel;
  wire   [3:0] comp_smpl;
  wire   [7:0] r_cvcwdat;
  wire   [7:0] r_sdischg;
  wire   [7:0] r_vcomp;
  wire   [7:0] r_idacsh;
  wire   [7:0] r_cvofsx;
  wire   [7:0] r_xtm;
  wire   [6:0] bist_r_ctl;
  wire   [1:0] regx_hitbst;
  wire   [7:0] bist_r_dat;
  wire   [1:0] regx_wrpwm;
  wire   [15:0] r_pwm;
  wire   [1:0] r_sap;
  wire   [3:0] lt_gpi;
  wire   [6:0] r_do_ts;
  wire   [3:0] r_dpdo_sel;
  wire   [3:0] r_dndo_sel;
  wire   [4:0] di_aswk;
  wire   [15:8] r_xana;
  wire   [4:0] di_xanav;
  wire   [7:0] r_aopt;
  wire   [6:0] di_gpio;
  wire   [7:6] do_opt;
  wire   [1:0] pwm_o;
  wire   [15:0] d_dodat;
  wire   [3:0] r_lt_gpi;
  tri   [7:0] SRAM_RDAT;

  CKBUFX1 U0_ASWCLK_BUF_0_ ( .A(aswclk_ps[0]), .Y(aswclk_ps[1]) );
  CKBUFX1 U0_ASWCLK_BUF_1_ ( .A(aswclk_ps[1]), .Y(aswclk_ps[2]) );
  CKBUFX1 U0_ASWCLK_BUF_2_ ( .A(aswclk_ps[2]), .Y(aswclk_ps[3]) );
  CKBUFX1 U0_ASWCLK_BUF_3_ ( .A(aswclk_ps[3]), .Y(aswclk_ps[4]) );
  CKBUFX1 U0_ASWCLK_BUF_4_ ( .A(aswclk_ps[4]), .Y(aswclk_ps[5]) );
  CKBUFX1 U0_ASWCLK_BUF_5_ ( .A(aswclk_ps[5]), .Y(aswclk_ps[6]) );
  CKBUFX1 U0_ASWCLK_BUF_6_ ( .A(aswclk_ps[6]), .Y(aswclk_ps[7]) );
  CKBUFX1 U0_ASWCLK_BUF_7_ ( .A(aswclk_ps[7]), .Y(aswclk_ps[8]) );
  CKBUFX1 U0_ASWCLK_BUF_8_ ( .A(aswclk_ps[8]), .Y(aswclk_ps[9]) );
  CKBUFX1 U0_ASWCLK_BUF_9_ ( .A(aswclk_ps[9]), .Y(aswclk) );
  CKBUFX1 U0_DETCLK_BUF_0_ ( .A(detclk_ps[0]), .Y(detclk_ps[1]) );
  CKBUFX1 U0_DETCLK_BUF_1_ ( .A(detclk_ps[1]), .Y(detclk_ps[2]) );
  CKBUFX1 U0_DETCLK_BUF_2_ ( .A(detclk_ps[2]), .Y(detclk_ps[3]) );
  CKBUFX1 U0_DETCLK_BUF_3_ ( .A(detclk_ps[3]), .Y(detclk_ps[4]) );
  CKBUFX1 U0_DETCLK_BUF_4_ ( .A(detclk_ps[4]), .Y(detclk_ps[5]) );
  CKBUFX1 U0_DETCLK_BUF_5_ ( .A(detclk_ps[5]), .Y(detclk_ps[6]) );
  CKBUFX1 U0_DETCLK_BUF_6_ ( .A(detclk_ps[6]), .Y(detclk_ps[7]) );
  CKBUFX1 U0_DETCLK_BUF_7_ ( .A(detclk_ps[7]), .Y(detclk_ps[8]) );
  CKBUFX1 U0_DETCLK_BUF_8_ ( .A(detclk_ps[8]), .Y(detclk_ps[9]) );
  CKBUFX1 U0_DETCLK_BUF_9_ ( .A(detclk_ps[9]), .Y(detclk) );
  AND2X1 U0_SCAN_EN ( .A(DI_GPIO[2]), .B(n72), .Y() );
  CKMUX2X1 U0_CLK_MUX ( .D0(i_clk), .D1(DI_GPIO[4]), .S(tclk_sel), .Y(s_clk)
         );
  CKMUX2X1 U0_DCLKMUX ( .D0(RD_DET), .D1(DI_GPIO[4]), .S(tclk_sel), .Y(
        detclk_ps[0]) );
  CKMUX2X1 U0_ACLKMUX ( .D0(aswkup), .D1(DI_GPIO[4]), .S(tclk_sel), .Y(
        aswclk_ps[0]) );
  CKBUFX1 U0_MCK_BUF ( .A(i_clk), .Y(x_clk) );
  CKBUFX1 U0_TCK_BUF ( .A(DI_GPIO[4]), .Y(t_di_gpio4) );
  CLKDLX1 U0_MCLK_ICG ( .CK(s_clk), .E(n573), .SE(n73), .ECK(g_clk) );
  CLKDLX1 U0_SRAM_ICG ( .CK(g_clk), .E(sram_en), .SE(n73), .ECK(SRAM_CLK) );
  INVX1 U0_REVIDZ_0_ ( .A(1'b1), .Y(REVID[0]) );
  INVX1 U0_REVIDZ_1_ ( .A(1'b1), .Y(REVID[1]) );
  INVX1 U0_REVIDZ_2_ ( .A(1'b1), .Y(REVID[2]) );
  INVX1 U0_REVIDZ_3_ ( .A(1'b1), .Y(REVID[3]) );
  INVX1 U0_REVIDZ_4_ ( .A(1'b0), .Y(REVID[4]) );
  INVX1 U0_REVIDZ_5_ ( .A(1'b0), .Y(REVID[5]) );
  INVX1 U0_REVIDZ_6_ ( .A(1'b1), .Y(REVID[6]) );
  mpb_a0 u0_mpb ( .i_rd({prl_cany0r, n77}), .i_wr({prl_cany0w, i2c_ev_3}), 
        .wdat0(sse_wdat), .wdat1(prx_fifowdat), .addr0(sse_adr), .addr1(
        prl_cany0adr), .r_i2c_attr(r_i2c_attr), .esfrm_oe(esfrm_oe), 
        .esfrm_we(esfrm_we), .sfrack(sfrack), .esfrm_wdat(esfrm_wdat), 
        .esfrm_adr(esfrm_adr), .mcu_esfr_rdat(mcu_esfrrdat), .delay_rdat(
        delay_inst), .delay_rrdy(ictlr_psrack), .esfrm_rrdy(esfrm_rrdy), 
        .esfrm_rdat(esfrm_rdat), .channel_sel(1'b0), .r_pg0_sel(r_pg0_sel), 
        .dma_w(1'b0), .dma_r(1'b0), .dma_addr({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .dma_wdat({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .dma_ack(), .memaddr(memaddr), 
        .memaddr_c({memaddr_c[15:5], n23, memaddr_c[3], n24, memaddr_c[1:0]}), 
        .memwr(memwr), .memrd(memrd), .memrd_c(memrd_c), .cpurst(o_cpurst), 
        .memdatao(memdatao), .memack(memack), .hit_xd(hit_xd), .hit_xr(hit_xr), 
        .hit_ps(hit_ps), .hit_ps_c(hit_ps_c), .idat_r(mcu_ram_r), .idat_w(
        mcu_ram_w), .idat_adr(idat_adr), .idat_wdat(idat_wdat), .iram_ce(
        iram_ce), .xram_ce(xram_ce), .regx_re(regx_re), .iram_we(iram_we), 
        .xram_we(xram_we), .regx_we(regx_we), .iram_a(iram_a), .xram_a(xram_a), 
        .iram_d(iram_d), .xram_d(xram_d), .iram_rdat({n136, n138, n140, n142, 
        n145, n147, sram_rdat}), .xram_rdat({n136, n138, n140, n142, n145, 
        n147, sram_rdat}), .regx_rdat(regx_rdat), .bist_en(n9), .bist_wr(
        bist_wr), .bist_adr(bist_adr), .bist_wdat(bist_wdat), .bist_xram(1'b0), 
        .mclk(g_clk), .srstz(n51) );
  mcu51_a0 u0_mcu ( .bclki2c(r_bclk_sel), .pc_ini({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .slp2wakeup(1'b0), .r_hold_mcu(r_hold_mcu), .wdt_slow(1'b0), .wdtov({
        SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2}), .mdubsy(), .cs_run(), 
        .t0_intr(t0_intr), .clki2c(g_clk), .clkmdu(g_clk), .clkur0(g_clk), 
        .clktm0(g_clk), .clktm1(g_clk), .clkwdt(g_clk), .i2c_autoack(1'b0), 
        .i2c_con_ens1(), .clkcpu(g_clk), .clkper(g_clk), .reset(n53), .ro(
        o_cpurst), .port0i({n587, di_gpio[6:4], n134, di_gpio[2:0]}), 
        .exint_9(fcp_intr), .exint({exint[7:4], n31, n30, exint[1:0]}), 
        .clkcpuen(), .clkperen(), .port0o({SYNOPSYS_UNCONNECTED_3, do_p0}), 
        .port0ff(ff_p0), .rxd0o(do_opt[7]), .txd0(do_opt[6]), .rxd0i(dpdm_urx), 
        .rxd0oe(s0_rxdoe), .scli(n505), .sdai(n507), .sclo(mcuo_scl), .sdao(
        mcuo_sda), .waitstaten(), .mempsack(mempsack), .memack(memack), 
        .memdatai(memdatai), .memdatao(memdatao), .memaddr(memaddr), .mempswr(
        mempswr), .mempsrd(mempsrd), .memwr(memwr), .memrd(memrd), 
        .memdatao_comb({SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5, 
        SYNOPSYS_UNCONNECTED_6, SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8, 
        SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10, 
        SYNOPSYS_UNCONNECTED_11}), .memaddr_comb(memaddr_c), .mempswr_comb(), 
        .mempsrd_comb(mempsrd_c), .memwr_comb(), .memrd_comb(memrd_c), 
        .ramdatai({n136, n138, n140, n142, n145, n147, sram_rdat}), .ramdatao(
        idat_wdat), .ramaddr(idat_adr), .ramwe(mcu_ram_w), .ramoe(mcu_ram_r), 
        .dbgpo({SYNOPSYS_UNCONNECTED_12, SYNOPSYS_UNCONNECTED_13, 
        SYNOPSYS_UNCONNECTED_14, SYNOPSYS_UNCONNECTED_15, 
        SYNOPSYS_UNCONNECTED_16, SYNOPSYS_UNCONNECTED_17, 
        SYNOPSYS_UNCONNECTED_18, SYNOPSYS_UNCONNECTED_19, 
        SYNOPSYS_UNCONNECTED_20, mcu_dbgpo, mcu_pc}), .sfrack(sfrack), 
        .sfrdatai(sfr_rdat), .sfrdatao(sfr_wdat), .sfraddr(sfr_adr), .sfrwe(
        sfr_w), .sfroe(sfr_r), .esfrm_wrdata(esfrm_wdat), .esfrm_addr(
        esfrm_adr), .esfrm_we(esfrm_we), .esfrm_oe(esfrm_oe), .esfrm_rddata(
        mcu_esfrrdat) );
  ictlr_a0 u0_ictlr ( .bkpt_ena(bkpt_ena), .bkpt_pc(bkpt_pc), .memaddr_c({
        memaddr_c[14:5], n23, memaddr_c[3], n24, n27, n26}), .memaddr(
        memaddr[14:0]), .mcu_psr_c(mempsrd_c), .mcu_psw(mempswr), .hit_ps_c(
        hit_ps_c), .hit_ps(hit_ps), .mempsack(ictlr_psack), .memdatao(memdatao), .o_set_hold(set_hold), .o_bkp_hold(bkpt_hold), .o_ofs_inc(ictlr_inc), 
        .o_inst(ictlr_inst), .d_inst(delay_inst), .sfr_psrack(ictlr_psrack), 
        .sfr_psofs(r_inst_ofs), .sfr_psr(r_psrd), .sfr_psw(r_pswr), .dw_rst(
        prl_c0set), .dw_ena(prl_cany0), .sfr_wdat({sfr_wdat[7], n47, n45, n42, 
        sfr_wdat[3:2], n35, n32}), .pmem_pgm(pmem_pgm), .pmem_re(pmem_re), 
        .pmem_csb(pmem_csb), .pmem_clk(pmem_clk), .pmem_a(PMEM_A), .pmem_q0(
        pmem_q0), .pmem_q1(pmem_q1), .pmem_twlb(pmem_twlb), .wd_twlb(wd_twlb), 
        .we_twlb(we_twlb), .pwrdn_rst(pwrdn_rst), .r_pwdn_en(r_otp_pwdn_en), 
        .r_multi(r_otp_wpls), .r_hold_mcu(r_hold_mcu), .clk(g_clk), .srst(
        o_cpurst) );
  regbank_a0 u0_regbank ( .srci({di_pro[5], n580, n581, n582, n583, di_pro[0]}), .dm_fault(di_aswk[3]), .cc1_di(n586), .cc2_di(n585), .di_rd_det(n122), 
        .di_stbovp(di_aswk[1]), .i_tmrf(t0_intr), .i_vcbyval(r_xtm[4]), 
        .dnchk_en(o_dodat5_2_), .r_pwrv_upd(r_pwrv_upd), .aswkup(aswkup), 
        .ps_pwrdn(ps_pwrdn), .r_sleep(r_sleep), .r_pwrdn(r_pwrdn), 
        .r_ocdrv_enz(r_ocdrv_enz), .r_osc_stop(r_osc_stop), .r_osc_lo(
        o_dodat0_15_), .r_osc_gate(r_osc_gate), .r_fw_pwrv(r_fw_pwrv), 
        .r_cvcwr(r_cvcwr[1:0]), .r_cvofs(r_cvofs), .r_otpi_gate(r_otpi_gate), 
        .r_pwrctl(r_pwrctl), .r_pwr_i(DO_PWR_I), .r_cvctl(r_cvctl), .r_srcctl(
        r_srcctl), .r_dpdmctl(r_dpdmctl), .r_ccrx({r_sqlch, 
        SYNOPSYS_UNCONNECTED_21, SYNOPSYS_UNCONNECTED_22, r_ccrx, r_rxdb_opt}), 
        .r_cctrx(r_cctrx), .r_ccctl(r_ccctl), .r_fcpwr(r_fcpwr), .r_fcpre(
        r_fcpre), .fcp_r_dat(fcp_r_dat), .fcp_r_sta(fcp_r_sta), .fcp_r_msk(
        fcp_r_msk), .fcp_r_ctl(fcp_r_ctl), .fcp_r_crc(fcp_r_crc), .fcp_r_acc(
        fcp_r_acc), .fcp_r_tui(fcp_r_tui), .r_accctl(r_accctl), .r_bclk_sel(
        r_bclk_sel), .r_dacwr(sfr_dacwr), .r_dac_en(r_dac_en[7:0]), .r_sar_en(
        r_sar_en[7:0]), .r_adofs({r_adofs[7], n14, n16, n15, n19, n17, n18, 
        r_adofs[0]}), .r_isofs(r_isofs), .x_daclsb(x_daclsb), .r_comp_opt({
        r_comp_opt, SYNOPSYS_UNCONNECTED_23, SYNOPSYS_UNCONNECTED_24, 
        SYNOPSYS_UNCONNECTED_25, SYNOPSYS_UNCONNECTED_26, 
        SYNOPSYS_UNCONNECTED_27}), .dac_r_ctl(dac_r_ctl), .dac_r_comp(
        dac_r_comp[7:0]), .dac_r_cmpsta(dac_r_cmpsta), .dac_r_vs(
        dac_r_vs[63:0]), .REVID(REVID), .atpg_en(n72), .sfr_r(sfr_r), .sfr_w(
        sfr_w), .set_hold(set_hold), .bkpt_hold(bkpt_hold), .cpurst(o_cpurst), 
        .sfr_addr({1'b1, sfr_adr}), .sfr_wdat({n49, n47, n44, n41, n39, n37, 
        n34, n28}), .sfr_rdat(sfr_rdat), .ff_p0(ff_p0), .di_p0({n587, 
        di_gpio[6:4], n134, di_gpio[2:0]}), .ictlr_idle(pmem_csb), .ictlr_inc(
        ictlr_inc), .r_inst_ofs(r_inst_ofs), .r_psrd(r_psrd), .r_pswr(r_pswr), 
        .r_fortxdat(r_fortxdat), .r_fortxrdy(r_fortxrdy), .r_fortxen(r_fortxen), .r_ana_tm(r_ana_tm), .r_gpio_tm(r_gpio_tm), .r_gpio_ie(r_gpio_ie), 
        .r_gpio_oe(r_gpio_oe), .r_gpio_pu(r_pu_gpio), .r_gpio_pd(r_pd_gpio), 
        .r_gpio_s0({N269, N268, N267}), .r_gpio_s1({N266, N265, N264}), 
        .r_gpio_s2({N263, N262, N261}), .r_gpio_s3({N260, N259, N258}), 
        .r_regtrm(r_regtrm), .i_pc(mcu_pc), .i_goidle(pid_goidle), .i_gobusy(
        pid_gobusy), .i_i2c_idle(sse_idle), .bus_idle(bus_idle), .i2c_stretch(
        hwi2c_stretch), .i_i2c_rwbuf(sse_wdat), .i_i2c_ltbuf(i2c_ltbuf), 
        .i_i2c_ofs(i2c_lt_ofs), .o_intr({exint[6], sfr_intr, exint[5:4]}), 
        .r_auto_gdcrc(r_auto_gdcrc), .r_exist1st(r_exist1st), .r_ordrs4(
        r_ordrs4), .r_fifopsh(r_fifopsh), .r_fifopop(r_fifopop), .r_unlock(
        r_unlock), .r_first(r_first), .r_last(r_last), .r_fiforst(r_fiforst), 
        .r_set_cpmsgid(r_set_cpmsgid), .r_txendk(r_txendk), .r_txnumk(r_txnumk), .r_txshrt(r_txshrt), .r_auto_discard(r_auto_discard), .r_hold_mcu(r_hold_mcu), .r_txauto(r_txauto), .r_rxords_ena(r_rxords_ena), .r_spec(r_spec), 
        .r_dat_spec(r_dat_spec), .r_dat_portrole(r_dat_portrole), 
        .r_dat_datarole(r_dat_datarole), .r_discard(r_discard), .r_pshords(
        r_pshords), .r_pg0_sel(r_pg0_sel), .r_strtch(r_strtch), .r_i2c_attr(
        r_i2c_attr), .r_i2c_ninc(r_i2c_ninc), .r_hwi2c_en(), .r_i2c_fwnak(
        r_i2c_fwnak), .r_i2c_fwack(r_i2c_fwack), .r_i2c_deva(r_i2c_deva), 
        .i2c_ev({n77, i2c_ev_6_, slvo_ev[3:2], i2c_ev_3, i2c_ev_2, 
        slvo_ev[1:0]}), .prl_c0set(prl_c0set), .prl_cany0(prl_cany0), 
        .prl_discard(prl_discard), .prl_GCTxDone(prl_GCTxDone), .prl_cpmsgid(
        prl_cpmsgid), .pff_ack(pff_ack), .prx_rst(prx_rst), .pff_obsd(pff_obsd), .pff_full(pff_full), .pff_empty(pff_empty), .ptx_ack(ptx_ack), .pff_ptr(
        pff_ptr), .prx_adpn(prx_adpn), .pff_rdat(pff_rdat), .pff_rxpart(
        pff_rxpart), .prx_rcvinf(prx_rcvinf), .ptx_fsm(ptx_fsm), .prx_fsm(
        prx_fsm), .prl_fsm(prl_fsm), .prx_setsta(prx_setsta), .clk_1500k(
        clk_1500k), .clk_500k(clk_500k), .clk_500(clk_500), .clk(g_clk), 
        .xrstz(i_rstz), .xclk(s_clk), .dbgpo({SYNOPSYS_UNCONNECTED_28, 
        SYNOPSYS_UNCONNECTED_29, SYNOPSYS_UNCONNECTED_30, 
        SYNOPSYS_UNCONNECTED_31, SYNOPSYS_UNCONNECTED_32, 
        SYNOPSYS_UNCONNECTED_33, SYNOPSYS_UNCONNECTED_34, 
        SYNOPSYS_UNCONNECTED_35, SYNOPSYS_UNCONNECTED_36, 
        SYNOPSYS_UNCONNECTED_37, SYNOPSYS_UNCONNECTED_38, 
        SYNOPSYS_UNCONNECTED_39, SYNOPSYS_UNCONNECTED_40, 
        SYNOPSYS_UNCONNECTED_41, SYNOPSYS_UNCONNECTED_42, 
        SYNOPSYS_UNCONNECTED_43, SYNOPSYS_UNCONNECTED_44, 
        SYNOPSYS_UNCONNECTED_45, SYNOPSYS_UNCONNECTED_46, 
        SYNOPSYS_UNCONNECTED_47, SYNOPSYS_UNCONNECTED_48, 
        SYNOPSYS_UNCONNECTED_49, SYNOPSYS_UNCONNECTED_50, 
        SYNOPSYS_UNCONNECTED_51, SYNOPSYS_UNCONNECTED_52, 
        SYNOPSYS_UNCONNECTED_53, SYNOPSYS_UNCONNECTED_54, 
        SYNOPSYS_UNCONNECTED_55, SYNOPSYS_UNCONNECTED_56, 
        SYNOPSYS_UNCONNECTED_57, SYNOPSYS_UNCONNECTED_58, 
        SYNOPSYS_UNCONNECTED_59}), .srstz(srstz), .prstz(prstz) );
  i2cslv_a0 u0_i2cslv ( .i_sda(n506), .i_scl(n504), .o_sda(slvo_sda), .i_deva(
        r_i2c_deva), .i_inc(n29), .i_fwnak(r_i2c_fwnak), .i_fwack(r_i2c_fwack), 
        .o_we(i2c_ev_3), .o_re(slvo_re), .o_r_early(slvo_early), .o_idle(
        sse_idle), .o_dec(), .o_busev(slvo_ev), .o_ofs(sse_adr), .o_lt_ofs(
        i2c_lt_ofs), .o_wdat(sse_wdat), .o_lt_buf(i2c_ltbuf), .o_dbgpo({
        SYNOPSYS_UNCONNECTED_60, SYNOPSYS_UNCONNECTED_61, 
        SYNOPSYS_UNCONNECTED_62, SYNOPSYS_UNCONNECTED_63, 
        SYNOPSYS_UNCONNECTED_64, SYNOPSYS_UNCONNECTED_65, 
        SYNOPSYS_UNCONNECTED_66, SYNOPSYS_UNCONNECTED_67}), .i_rdat(esfrm_rdat), .i_rd_mem(sse_rdrdy), .i_clk(g_clk), .i_rstz(n52), .i_prefetch(sse_prefetch)
         );
  updphy_FF_DEPTH_NUM34_FF_DEPTH_NBT6 u0_updphy ( .i_cc(di_cc), .i_cc_49(n584), 
        .i_sqlch(n124), .r_sqlch(r_sqlch), .r_adprx_en(r_ccrx[3]), .r_adp2nd(
        r_ccrx[2]), .r_exist1st(r_exist1st), .r_ordrs4(r_ordrs4), .r_fifopsh(
        r_fifopsh), .r_fifopop(r_fifopop), .r_fiforst(r_fiforst), .r_unlock(
        r_unlock), .r_first(r_first), .r_last(r_last), .r_set_cpmsgid(
        r_set_cpmsgid), .r_rdy(upd_rdrdy), .r_wdat({n49, n47, n45, n42, 
        sfr_wdat[3], n37, n35, n32}), .r_rdat(esfrm_rdat), .r_txnumk(r_txnumk), 
        .r_txendk(r_txendk), .r_txshrt(r_txshrt), .r_auto_discard(
        r_auto_discard), .r_txauto(r_txauto), .r_rxords_ena(r_rxords_ena), 
        .r_spec(r_spec), .r_dat_spec(r_dat_spec), .r_auto_gdcrc(r_auto_gdcrc), 
        .r_rxdb_opt(r_rxdb_opt), .r_pshords(r_pshords), .r_dat_portrole(
        r_dat_portrole), .r_dat_datarole(r_dat_datarole), .r_discard(r_discard), .pid_goidle(pid_goidle), .pid_gobusy(pid_gobusy), .pff_ack(pff_ack), 
        .pff_rdat(pff_rdat), .pff_rxpart(pff_rxpart), .prx_rcvinf(prx_rcvinf), 
        .pff_obsd(pff_obsd), .pff_ptr(pff_ptr), .pff_empty(pff_empty), 
        .pff_full(pff_full), .ptx_ack(ptx_ack), .ptx_cc(ptx_cc), .ptx_oe(
        ptx_oe), .prx_setsta(prx_setsta), .prx_rst(prx_rst), .prl_c0set(
        prl_c0set), .prl_cany0(prl_cany0), .prl_cany0r(prl_cany0r), 
        .prl_cany0w(prl_cany0w), .prl_discard(prl_discard), .prl_GCTxDone(
        prl_GCTxDone), .prl_cany0adr(prl_cany0adr), .prl_cpmsgid(prl_cpmsgid), 
        .prx_fifowdat(prx_fifowdat), .ptx_fsm(ptx_fsm), .prl_fsm(prl_fsm), 
        .prx_fsm(prx_fsm), .prx_adpn(prx_adpn), .dbgpo({
        SYNOPSYS_UNCONNECTED_68, SYNOPSYS_UNCONNECTED_69, 
        SYNOPSYS_UNCONNECTED_70, SYNOPSYS_UNCONNECTED_71, 
        SYNOPSYS_UNCONNECTED_72, SYNOPSYS_UNCONNECTED_73, 
        SYNOPSYS_UNCONNECTED_74, SYNOPSYS_UNCONNECTED_75, 
        SYNOPSYS_UNCONNECTED_76, SYNOPSYS_UNCONNECTED_77, 
        SYNOPSYS_UNCONNECTED_78, SYNOPSYS_UNCONNECTED_79, 
        SYNOPSYS_UNCONNECTED_80, upd_dbgpo, SYNOPSYS_UNCONNECTED_81, 
        SYNOPSYS_UNCONNECTED_82, SYNOPSYS_UNCONNECTED_83, 
        SYNOPSYS_UNCONNECTED_84, SYNOPSYS_UNCONNECTED_85, 
        SYNOPSYS_UNCONNECTED_86, SYNOPSYS_UNCONNECTED_87, 
        SYNOPSYS_UNCONNECTED_88, SYNOPSYS_UNCONNECTED_89, 
        SYNOPSYS_UNCONNECTED_90, SYNOPSYS_UNCONNECTED_91, 
        SYNOPSYS_UNCONNECTED_92, SYNOPSYS_UNCONNECTED_93, 
        SYNOPSYS_UNCONNECTED_94, SYNOPSYS_UNCONNECTED_95, 
        SYNOPSYS_UNCONNECTED_96, SYNOPSYS_UNCONNECTED_97}), .clk(g_clk), 
        .srstz(prstz) );
  dacmux_a0 u0_dacmux ( .clk(g_clk), .srstz(n51), .i_comp(n587), .r_comp_opt(
        r_comp_opt), .r_wdat(r_dacwdat), .r_adofs(r_adofs), .r_isofs(r_isofs), 
        .r_wr({r_dacwr, sfr_dacwr[14:8]}), .dacv_wr({wr_dacv[17:16], n25, 
        wr_dacv[14:8], sfr_dacwr[7:0]}), .o_dacv(dac_r_vs), .o_shrst(sh_rst), 
        .o_hold(sh_hold), .o_dac1(DAC1_V), .o_daci_sel(dacmux_sel), .o_dat(
        dac_r_comp), .r_dac_en(r_dac_en), .r_sar_en(r_sar_en), .o_dactl(
        dac_r_ctl), .o_cmpsta(dac_r_cmpsta), .x_daclsb(x_daclsb), .o_intr(
        exint[7]), .o_smpl({SYNOPSYS_UNCONNECTED_98, comp_smpl}) );
  fcp_a0 u0_fcp ( .dp_comp(dp_comp), .dm_comp(dm_comp), .id_comp(1'b0), .intr(
        fcp_intr), .tx_en(fcp_oe), .tx_dat(fcp_do), .r_dat(fcp_r_dat), .r_sta(
        fcp_r_sta), .r_ctl(fcp_r_ctl), .r_msk(fcp_r_msk), .r_crc(fcp_r_crc), 
        .r_acc(fcp_r_acc), .r_dpdmsta(r_accctl), .r_wdat({n49, n47, n45, n42, 
        n39, n37, n35, n32}), .r_wr(r_fcpwr), .r_re(r_fcpre), .clk(g_clk), 
        .srstz(n52), .r_tui(fcp_r_tui) );
  cvctl_a0 u0_cvctl ( .r_cvcwr(r_cvcwr), .wdat(r_cvcwdat), .r_sdischg(
        r_sdischg), .r_vcomp(r_vcomp), .r_idacsh(r_idacsh), .r_cvofsx(r_cvofsx), .r_cvofs(r_cvofs), .sdischg_duty(sdischg_duty), .r_hlsb_en(r_pwrctl[4]), 
        .r_hlsb_sel(r_pwrctl[5]), .r_hlsb_freq(r_xtm[5]), .r_hlsb_duty(
        r_xtm[6]), .r_fw_pwrv(r_fw_pwrv), .r_dac0(DO_DAC0), .r_dac3(DAC3_V), 
        .clk_100k(clk_100k), .clk(g_clk), .srstz(n52) );
  regx_a0 u0_regx ( .regx_r(regx_re), .regx_w(regx_we), .di_drposc(di_aswk[0]), 
        .di_imposc(di_aswk[4]), .di_rd_det(n122), .di_stbovp(di_aswk[1]), 
        .clk_500k(clk_500k), .r_imp_osc(r_imp_osc), .regx_addr({xram_a[6:5], 
        n1, xram_a[3:0]}), .regx_wdat(xram_d), .regx_rdat(regx_rdat), 
        .regx_hitbst(regx_hitbst), .regx_wrpwm(regx_wrpwm), .regx_wrcvc({
        r_cvcwr[2], r_cvcwr[5:3]}), .r_sdischg(r_sdischg), .r_bistctl(
        bist_r_ctl), .r_bistdat(bist_r_dat), .r_vcomp(r_vcomp), .r_idacsh(
        r_idacsh), .r_cvofsx(r_cvofsx), .r_pwm(r_pwm), .regx_wrdac({
        wr_dacv[17:16], r_dacwr[10:9], wr_dacv[15:8], r_dacwr[8:7]}), 
        .dac_r_vs(dac_r_vs[143:64]), .dac_comp(dac_r_comp[17:8]), .r_dac_en(
        r_dac_en[17:8]), .r_sar_en(r_sar_en[17:8]), .r_aopt(r_aopt), .r_xtm(
        r_xtm), .r_adummyi(DUMMY_IN), .r_bck0(BCK_REGX[7:0]), .r_bck1(
        BCK_REGX[15:8]), .r_i2crout({r_i2crout, r_i2cmcu_route, r_i2cslv_route}), .r_xana({r_xana_23, SYNOPSYS_UNCONNECTED_99, SYNOPSYS_UNCONNECTED_100, 
        SYNOPSYS_UNCONNECTED_101, r_xana_19, r_xana_18, OCP_SEL, PWREN_HOLD, 
        r_xana, ANA_REGX[7:0]}), .di_xana(di_xanav), .lt_gpi(lt_gpi), .di_tst(
        di_tst), .bkpt_pc(bkpt_pc), .bkpt_ena(bkpt_ena), .we_twlb(we_twlb), 
        .r_vpp_en(r_vpp_en), .r_vpp0v_en(r_vpp0v_en), .r_otp_pwdn_en(
        r_otp_pwdn_en), .r_otp_wpls(r_otp_wpls), .wd_twlb(wd_twlb), .r_sap(
        r_sap), .r_twlb(pmem_twlb), .upd_pwrv(r_pwrv_upd), .ramacc(ramacc), 
        .sse_idle(sse_idle), .bus_idle(bus_idle), .r_do_ts(r_do_ts), 
        .r_dpdo_sel(r_dpdo_sel), .r_dndo_sel(r_dndo_sel), .di_ts(di_ts), 
        .detclk(detclk), .aswclk(aswclk), .atpg_en(n72), .di_aswk({
        di_aswk[4:3], n122, di_aswk[1:0]}), .clk(g_clk), .rrstz(srstz) );
  srambist_a0 u0_srambist ( .clk(g_clk), .srstz(n52), .reg_hit(regx_hitbst), 
        .reg_w(regx_we), .reg_r(regx_re), .reg_wdat(xram_d), .iram_rdat({n136, 
        n138, n140, n142, n145, n147, sram_rdat}), .xram_rdat({n136, n138, 
        n140, n142, n145, n147, sram_rdat}), .bist_en(bist_en), .bist_xram(), 
        .bist_wr(bist_wr), .bist_adr(bist_adr), .bist_wdat(bist_wdat), 
        .o_bistctl(bist_r_ctl), .o_bistdat(bist_r_dat) );
  divclk_a0 u0_divclk ( .mclk(g_clk), .srstz(n52), .atpg_en(n54), .clk_1500k(
        clk_1500k), .clk_500k(clk_500k), .clk_100k(clk_100k), .clk_50k(clk_50k), .clk_500(clk_500), .divff_8(divff_8), .divff_5(divff_5) );
  glpwm_a0_0 u0_pwm_0_ ( .clk(g_clk), .rstz(n52), .clk_base(clk_50k), .we(
        regx_wrpwm[0]), .wdat(xram_d), .r_pwm(r_pwm[7:0]), .pwm_o(pwm_o[0]) );
  glpwm_a0_1 u0_pwm_1_ ( .clk(g_clk), .rstz(n51), .clk_base(clk_50k), .we(
        regx_wrpwm[1]), .wdat(xram_d), .r_pwm(r_pwm[15:8]), .pwm_o(pwm_o[1])
         );
  SNPS_CLOCK_GATE_HIGH_core_a0 clk_gate_d_dodat_reg ( .CLK(g_clk), .EN(N570), 
        .ENCLK(net8831), .TE(1'b0) );
  DLNQX1 r_lt_gpi_reg_1_ ( .D(DI_GPIO[2]), .XG(i_rstz), .Q(r_lt_gpi[1]) );
  DLNQX1 r_lt_gpi_reg_0_ ( .D(DI_GPIO[3]), .XG(i_rstz), .Q(r_lt_gpi[0]) );
  DLNQX1 r_lt_gpi_reg_2_ ( .D(DI_GPIO[1]), .XG(i_rstz), .Q(r_lt_gpi[2]) );
  DLNQX1 r_lt_gpi_reg_3_ ( .D(DI_GPIO[0]), .XG(i_rstz), .Q(r_lt_gpi[3]) );
  DFFQX1 d_dodat_reg_11_ ( .D(N1483), .C(net8831), .Q(d_dodat[11]) );
  DFFQX1 d_dodat_reg_12_ ( .D(N574), .C(net8831), .Q(d_dodat[12]) );
  DFFQX1 d_dodat_reg_14_ ( .D(N572), .C(net8831), .Q(d_dodat[14]) );
  DFFQX1 d_dodat_reg_8_ ( .D(N1498), .C(net8831), .Q(d_dodat[8]) );
  DFFQX1 d_dodat_reg_10_ ( .D(N1488), .C(net8831), .Q(d_dodat[10]) );
  DFFQX1 d_dodat_reg_9_ ( .D(N1493), .C(net8831), .Q(d_dodat[9]) );
  DFFQX1 d_dodat_reg_15_ ( .D(N571), .C(net8831), .Q(d_dodat[15]) );
  DFFQX1 d_dodat_reg_13_ ( .D(N573), .C(net8831), .Q(d_dodat[13]) );
  DFFQX1 d_dodat_reg_4_ ( .D(N582), .C(net8831), .Q(d_dodat[4]) );
  DFFQX1 d_dodat_reg_1_ ( .D(N585), .C(net8831), .Q(d_dodat[1]) );
  DFFQX1 d_dodat_reg_0_ ( .D(N586), .C(net8831), .Q(d_dodat[0]) );
  DFFQX1 d_dodat_reg_3_ ( .D(N583), .C(net8831), .Q(d_dodat[3]) );
  DFFQX1 d_dodat_reg_5_ ( .D(N581), .C(net8831), .Q(d_dodat[5]) );
  DFFQX1 d_dodat_reg_6_ ( .D(N580), .C(net8831), .Q(d_dodat[6]) );
  DFFQX1 d_dodat_reg_2_ ( .D(N584), .C(net8831), .Q(d_dodat[2]) );
  DFFQX1 d_dodat_reg_7_ ( .D(N579), .C(net8831), .Q(d_dodat[7]) );
  BUFX1 U3 ( .A(xram_a[4]), .Y(n1) );
  BUFXL U4 ( .A(n105), .Y(n2) );
  OA21X1 U5 ( .B(hit_xd), .C(hit_xr), .A(memrd), .Y(n3) );
  BUFX2 U6 ( .A(xram_ce), .Y(n4) );
  INVXL U7 ( .A(n3), .Y(n5) );
  INVXL U8 ( .A(n3), .Y(n6) );
  INVXL U9 ( .A(n630), .Y(n7) );
  INVX24 U10 ( .A(n7), .Y(PMEM_PGM) );
  NOR21XL U11 ( .B(pmem_pgm), .A(n73), .Y(n630) );
  BUFX3 U12 ( .A(bist_en), .Y(n9) );
  BUFX3 U13 ( .A(iram_ce), .Y(n10) );
  INVX1 U14 ( .A(n500), .Y(n11) );
  BUFX3 U15 ( .A(n627), .Y(PMEM_TWLB[0]) );
  NOR21XL U16 ( .B(pmem_twlb[0]), .A(n89), .Y(n627) );
  BUFX3 U17 ( .A(n499), .Y(n13) );
  BUFX3 U18 ( .A(r_adofs[6]), .Y(n14) );
  BUFX3 U19 ( .A(r_adofs[4]), .Y(n15) );
  BUFX3 U20 ( .A(r_adofs[5]), .Y(n16) );
  BUFX3 U21 ( .A(r_adofs[2]), .Y(n17) );
  BUFX3 U22 ( .A(r_adofs[1]), .Y(n18) );
  BUFX3 U23 ( .A(r_adofs[3]), .Y(n19) );
  BUFX3 U24 ( .A(n626), .Y(PMEM_TWLB[1]) );
  NOR21XL U25 ( .B(pmem_twlb[1]), .A(n89), .Y(n626) );
  BUFX4 U26 ( .A(n629), .Y(PMEM_SAP[0]) );
  NOR21XL U27 ( .B(r_sap[0]), .A(n90), .Y(n629) );
  BUFX4 U28 ( .A(n628), .Y(PMEM_SAP[1]) );
  NOR21XL U29 ( .B(r_sap[1]), .A(n91), .Y(n628) );
  OR2X2 U30 ( .A(r_dacwr[10]), .B(r_dacwr[9]), .Y(n102) );
  NOR3XL U31 ( .A(r_cvcwr[5]), .B(r_cvcwr[4]), .C(r_cvcwr[3]), .Y(n167) );
  AO22XL U32 ( .A(xram_a[0]), .B(xram_ce), .C(iram_a[0]), .D(iram_ce), .Y(
        SRAM_A[0]) );
  AOI221XL U33 ( .A(N634), .B(n499), .C(N600), .D(n569), .E(n600), .Y(n455) );
  AOI221XL U34 ( .A(N629), .B(n499), .C(N596), .D(n11), .E(n576), .Y(n353) );
  AOI221XL U35 ( .A(N644), .B(n499), .C(N610), .D(n569), .E(n595), .Y(n473) );
  AOI221XL U36 ( .A(N632), .B(n499), .C(N598), .D(n569), .E(n598), .Y(n456) );
  AOI221XL U37 ( .A(N637), .B(n499), .C(N603), .D(n569), .E(n590), .Y(n458) );
  AOI221XL U38 ( .A(N638), .B(n499), .C(N604), .D(n569), .E(n596), .Y(n471) );
  AOI221XL U39 ( .A(N633), .B(n499), .C(N599), .D(n11), .E(n592), .Y(n467) );
  AOI221XL U40 ( .A(N631), .B(n13), .C(N597), .D(n569), .E(n599), .Y(n481) );
  AOI221XL U41 ( .A(N640), .B(n13), .C(N606), .D(n11), .E(n589), .Y(n497) );
  AOI221XL U42 ( .A(N642), .B(n13), .C(N608), .D(n569), .E(n588), .Y(n482) );
  AOI221XL U43 ( .A(N641), .B(n13), .C(N607), .D(n11), .E(n594), .Y(n495) );
  AOI222XL U44 ( .A(N643), .B(n499), .C(N609), .D(n11), .E(d_dodat[14]), .F(
        n72), .Y(n472) );
  AOI22AXL U45 ( .A(r_fortxrdy), .B(r_fortxdat), .D(r_fortxrdy), .C(ptx_cc), 
        .Y(n321) );
  NOR21XL U46 ( .B(r_aopt[1]), .A(n62), .Y(ANAOPT[1]) );
  NOR21XL U47 ( .B(r_aopt[4]), .A(n62), .Y(ANAOPT[4]) );
  NOR21XL U48 ( .B(r_xana[8]), .A(n63), .Y(ANA_REGX[8]) );
  NOR21XL U49 ( .B(r_xana[9]), .A(n66), .Y(ANA_REGX[9]) );
  NOR21XL U50 ( .B(r_ccctl[1]), .A(n63), .Y(DO_CCCTL[1]) );
  NOR21XL U51 ( .B(r_ccctl[2]), .A(n63), .Y(DO_CCCTL[2]) );
  NOR21XL U52 ( .B(r_ccctl[3]), .A(n63), .Y(DO_CCCTL[3]) );
  NOR21XL U53 ( .B(r_cvctl[3]), .A(n65), .Y(DO_CVCTL[3]) );
  NOR21XL U54 ( .B(r_cvctl[4]), .A(n65), .Y(DO_CVCTL[4]) );
  NOR21XL U55 ( .B(r_srcctl[6]), .A(n66), .Y(DO_SRCCTL[6]) );
  NOR21XL U56 ( .B(r_srcctl[7]), .A(n67), .Y(DO_SRCCTL[7]) );
  OR2X1 U57 ( .A(r_cvctl[1]), .B(n73), .Y(DO_CVCTL[1]) );
  OR2X1 U58 ( .A(r_cvctl[0]), .B(n72), .Y(DO_CVCTL[0]) );
  OR2X1 U59 ( .A(wr_dacv[10]), .B(wr_dacv[9]), .Y(n99) );
  INVX1 U60 ( .A(n167), .Y(n118) );
  INVX1 U61 ( .A(n449), .Y(n557) );
  INVX1 U62 ( .A(n80), .Y(n60) );
  INVX1 U63 ( .A(n92), .Y(n59) );
  INVX1 U64 ( .A(n79), .Y(n58) );
  INVX1 U65 ( .A(n76), .Y(n57) );
  INVX1 U66 ( .A(n78), .Y(n61) );
  INVX1 U67 ( .A(n79), .Y(n56) );
  INVX1 U68 ( .A(n80), .Y(n55) );
  INVX1 U69 ( .A(n93), .Y(n64) );
  INVX1 U70 ( .A(n85), .Y(n62) );
  INVX1 U71 ( .A(n84), .Y(n63) );
  INVX1 U72 ( .A(n76), .Y(n65) );
  INVX1 U73 ( .A(n78), .Y(n66) );
  INVX1 U74 ( .A(n75), .Y(n67) );
  INVX1 U75 ( .A(n81), .Y(n68) );
  INVX1 U76 ( .A(n79), .Y(n54) );
  INVX1 U77 ( .A(n92), .Y(n69) );
  INVX1 U78 ( .A(n78), .Y(n70) );
  INVX1 U79 ( .A(n74), .Y(n71) );
  INVX1 U80 ( .A(n74), .Y(n72) );
  INVX1 U81 ( .A(n75), .Y(n73) );
  NAND21X1 U82 ( .B(wr_dacv[17]), .A(n96), .Y(n103) );
  NAND21X1 U83 ( .B(wr_dacv[15]), .A(n95), .Y(n104) );
  BUFXL U84 ( .A(wr_dacv[15]), .Y(n25) );
  INVX1 U85 ( .A(wr_dacv[11]), .Y(n98) );
  INVX1 U86 ( .A(wr_dacv[14]), .Y(n95) );
  INVX1 U87 ( .A(n40), .Y(n39) );
  INVX1 U88 ( .A(wr_dacv[16]), .Y(n96) );
  INVX1 U89 ( .A(r_dacwr[8]), .Y(n97) );
  NAND2X1 U90 ( .A(n92), .B(sram_en), .Y(SRAM_CEB) );
  INVX1 U91 ( .A(n33), .Y(n32) );
  INVX1 U92 ( .A(n48), .Y(n47) );
  INVX1 U93 ( .A(n38), .Y(n37) );
  INVX1 U94 ( .A(n53), .Y(n51) );
  INVX1 U95 ( .A(n50), .Y(n49) );
  INVX1 U96 ( .A(n43), .Y(n41) );
  INVX1 U97 ( .A(n33), .Y(n28) );
  INVX1 U98 ( .A(n36), .Y(n34) );
  INVX1 U99 ( .A(n46), .Y(n44) );
  INVX1 U100 ( .A(n36), .Y(n35) );
  INVX1 U101 ( .A(n43), .Y(n42) );
  INVX1 U102 ( .A(n46), .Y(n45) );
  NOR2X1 U103 ( .A(n352), .B(n561), .Y(n449) );
  INVX1 U104 ( .A(n53), .Y(n52) );
  INVX1 U105 ( .A(n90), .Y(n86) );
  INVX1 U106 ( .A(n90), .Y(n75) );
  INVX1 U107 ( .A(n91), .Y(n74) );
  INVX1 U108 ( .A(atpg_en), .Y(n76) );
  INVX1 U109 ( .A(n89), .Y(n78) );
  INVX1 U110 ( .A(atpg_en), .Y(n79) );
  INVX1 U111 ( .A(n89), .Y(n88) );
  INVX1 U112 ( .A(n89), .Y(n87) );
  INVX1 U113 ( .A(n73), .Y(n80) );
  INVX1 U114 ( .A(n91), .Y(n81) );
  INVX1 U115 ( .A(n91), .Y(n82) );
  INVX1 U116 ( .A(n90), .Y(n85) );
  INVX1 U117 ( .A(n90), .Y(n84) );
  INVX1 U118 ( .A(n91), .Y(n83) );
  NOR2X1 U119 ( .A(n70), .B(n129), .Y(OSC_LOW) );
  INVX1 U120 ( .A(sfr_wdat[3]), .Y(n40) );
  XNOR2XL U121 ( .A(n248), .B(DO_GPIO[2]), .Y(n269) );
  INVX1 U122 ( .A(n248), .Y(SRAM_A[2]) );
  INVX1 U123 ( .A(n247), .Y(SRAM_A[4]) );
  XNOR2XL U124 ( .A(n246), .B(SRAM_D[1]), .Y(n284) );
  XNOR2XL U125 ( .A(n245), .B(SRAM_D[2]), .Y(n289) );
  OR2X1 U126 ( .A(xram_ce), .B(iram_ce), .Y(sram_en) );
  INVX1 U127 ( .A(n246), .Y(SRAM_A[5]) );
  INVX1 U128 ( .A(n245), .Y(SRAM_A[6]) );
  OAI22X1 U129 ( .A(n167), .B(n120), .C(n36), .D(n118), .Y(r_cvcwdat[1]) );
  OAI22X1 U130 ( .A(n167), .B(n121), .C(n38), .D(n118), .Y(r_cvcwdat[2]) );
  OAI22XL U131 ( .A(n167), .B(n123), .C(n40), .D(n118), .Y(r_cvcwdat[3]) );
  OAI22X1 U132 ( .A(n167), .B(n127), .C(n48), .D(n118), .Y(r_cvcwdat[6]) );
  OAI22X1 U133 ( .A(n167), .B(n128), .C(n50), .D(n118), .Y(r_cvcwdat[7]) );
  INVX1 U134 ( .A(n242), .Y(SRAM_D[5]) );
  INVX1 U135 ( .A(n243), .Y(SRAM_D[4]) );
  XNOR2XL U136 ( .A(DAC3_V[4]), .B(n244), .Y(n276) );
  INVX1 U137 ( .A(n244), .Y(SRAM_D[0]) );
  INVX1 U138 ( .A(srstz), .Y(n53) );
  INVX1 U139 ( .A(sfr_wdat[0]), .Y(n33) );
  INVX1 U140 ( .A(sfr_wdat[2]), .Y(n38) );
  INVX1 U141 ( .A(sfr_wdat[6]), .Y(n48) );
  INVX1 U142 ( .A(sfr_wdat[7]), .Y(n50) );
  INVX1 U143 ( .A(sfr_wdat[5]), .Y(n46) );
  INVX1 U144 ( .A(sfr_wdat[1]), .Y(n36) );
  INVX1 U145 ( .A(sfr_wdat[4]), .Y(n43) );
  INVX1 U146 ( .A(xram_we), .Y(n119) );
  OAI21X1 U147 ( .B(xram_we), .C(iram_we), .A(n79), .Y(SRAM_WEB) );
  OR2X1 U148 ( .A(iram_we), .B(xram_we), .Y(n319) );
  NAND21X1 U149 ( .B(n465), .A(n455), .Y(n494) );
  INVX1 U150 ( .A(n338), .Y(do_opt_0) );
  NAND4X1 U151 ( .A(n473), .B(n482), .C(n471), .D(n458), .Y(n488) );
  NAND2X1 U152 ( .A(n459), .B(n453), .Y(n464) );
  NAND4X1 U153 ( .A(n497), .B(n467), .C(n495), .D(n498), .Y(n352) );
  NOR4XL U154 ( .A(n494), .B(n464), .C(n448), .D(n488), .Y(n498) );
  NAND2X1 U155 ( .A(n456), .B(n481), .Y(n465) );
  INVX1 U156 ( .A(n353), .Y(n561) );
  NAND2X1 U157 ( .A(n353), .B(n557), .Y(n487) );
  XNOR2XL U158 ( .A(DAC3_V[0]), .B(n523), .Y(n260) );
  NAND21X1 U159 ( .B(n448), .A(n473), .Y(n478) );
  INVX1 U160 ( .A(n467), .Y(n567) );
  INVX1 U161 ( .A(n455), .Y(n556) );
  INVX1 U162 ( .A(n482), .Y(n565) );
  INVX1 U163 ( .A(n458), .Y(n563) );
  INVX1 U164 ( .A(n471), .Y(n564) );
  INVX1 U165 ( .A(n481), .Y(n558) );
  INVX1 U166 ( .A(s0_rxdoe), .Y(n570) );
  INVX1 U167 ( .A(n497), .Y(n568) );
  INVX1 U168 ( .A(n495), .Y(n560) );
  INVX1 U169 ( .A(n473), .Y(n566) );
  INVX1 U170 ( .A(n456), .Y(n559) );
  INVX1 U171 ( .A(o_dodat0_15_), .Y(n129) );
  INVX1 U172 ( .A(n381), .Y(n219) );
  NOR2X1 U173 ( .A(n155), .B(n150), .Y(n360) );
  NOR21XL U174 ( .B(r_osc_stop), .A(n89), .Y(OSC_STOP) );
  NAND2X1 U175 ( .A(n601), .B(n602), .Y(n621) );
  NAND2X1 U176 ( .A(n579), .B(n578), .Y(n611) );
  NAND2X1 U177 ( .A(n94), .B(n154), .Y(tclk_sel) );
  INVX1 U178 ( .A(n94), .Y(n89) );
  INVX1 U179 ( .A(n93), .Y(n91) );
  INVX1 U180 ( .A(n94), .Y(n90) );
  AOI21X1 U181 ( .B(n153), .C(n149), .A(n73), .Y(CCI2C_EN) );
  NOR2X1 U182 ( .A(n71), .B(n137), .Y(ANAOPT[3]) );
  NAND2X1 U183 ( .A(n554), .B(n74), .Y(OCDRV_ENZ) );
  NAND2X1 U184 ( .A(n525), .B(n75), .Y(SH_HOLD) );
  INVX1 U185 ( .A(n154), .Y(n576) );
  BUFXL U186 ( .A(memaddr_c[0]), .Y(n26) );
  NOR21XL U187 ( .B(n295), .A(n67), .Y(DO_TS[3]) );
  XNOR2XL U188 ( .A(DO_GPIO[4]), .B(n247), .Y(n278) );
  XNOR2XL U189 ( .A(n266), .B(n267), .Y(N584) );
  XNOR2XL U190 ( .A(DAC3_V[2]), .B(n268), .Y(n267) );
  XNOR2XL U191 ( .A(n269), .B(n137), .Y(n266) );
  XNOR2XL U192 ( .A(DO_PWR_I[2]), .B(n526), .Y(n268) );
  XNOR2XL U193 ( .A(n274), .B(n275), .Y(N582) );
  XNOR2XL U194 ( .A(n276), .B(n277), .Y(n275) );
  XNOR2XL U195 ( .A(n278), .B(n279), .Y(n274) );
  XNOR2XL U196 ( .A(dacmux_sel[4]), .B(DO_PWR_I[4]), .Y(n277) );
  AOI22X1 U197 ( .A(n493), .B(n560), .C(n494), .D(n124), .Y(n492) );
  NAND2X1 U198 ( .A(n574), .B(n575), .Y(n493) );
  AOI22X1 U199 ( .A(pmem_csb), .B(n560), .C(n565), .D(dm_comp), .Y(n474) );
  NAND4X1 U200 ( .A(n489), .B(n490), .C(n491), .D(n492), .Y(DO_GPIO[2]) );
  AOI22AXL U201 ( .A(n568), .B(n587), .D(n470), .C(r_osc_stop), .Y(n489) );
  AOI22AXL U202 ( .A(n567), .B(n586), .D(n459), .C(di_pro[5]), .Y(n490) );
  AOI22X1 U203 ( .A(mcu_dbgpo[20]), .B(n496), .C(N450), .D(n487), .Y(n491) );
  OAI211X1 U204 ( .C(n156), .D(n207), .A(n208), .B(n209), .Y(memdatai[7]) );
  AOI22X1 U205 ( .A(regx_rdat[7]), .B(n210), .C(ictlr_inst[7]), .D(n6), .Y(
        n209) );
  AOI22XL U206 ( .A(xram_a[6]), .B(xram_ce), .C(iram_a[6]), .D(iram_ce), .Y(
        n245) );
  AOI22X1 U207 ( .A(xram_a[5]), .B(xram_ce), .C(iram_a[5]), .D(iram_ce), .Y(
        n246) );
  AO22X1 U208 ( .A(xram_a[3]), .B(xram_ce), .C(iram_a[3]), .D(iram_ce), .Y(
        SRAM_A[3]) );
  XNOR2XL U209 ( .A(sram_en), .B(n249), .Y(n312) );
  XNOR2XL U210 ( .A(SRAM_D[3]), .B(SRAM_A[7]), .Y(n294) );
  XNOR2XL U211 ( .A(n270), .B(n271), .Y(N583) );
  XNOR2XL U212 ( .A(DAC3_V[3]), .B(n272), .Y(n271) );
  XNOR2XL U213 ( .A(CC1_DOB), .B(n273), .Y(n270) );
  XNOR2XL U214 ( .A(DO_PWR_I[3]), .B(n527), .Y(n272) );
  XNOR2XL U215 ( .A(DO_GPIO[3]), .B(SRAM_A[3]), .Y(n273) );
  XNOR2XL U216 ( .A(n285), .B(n286), .Y(N580) );
  XNOR2XL U217 ( .A(n287), .B(n288), .Y(n286) );
  XOR2X1 U218 ( .A(DO_GPIO[6]), .B(n289), .Y(n285) );
  XNOR2XL U219 ( .A(DO_DAC0[1]), .B(DAC1_V[0]), .Y(n287) );
  XNOR2XL U220 ( .A(n280), .B(n281), .Y(N581) );
  XNOR2XL U221 ( .A(n282), .B(n283), .Y(n281) );
  XNOR2XL U222 ( .A(n284), .B(DO_GPIO[5]), .Y(n280) );
  XNOR2XL U223 ( .A(DO_DAC0[0]), .B(DAC3_V[5]), .Y(n282) );
  XNOR2XL U224 ( .A(n290), .B(n291), .Y(N579) );
  XNOR2XL U225 ( .A(n292), .B(n293), .Y(n291) );
  XNOR2XL U226 ( .A(n294), .B(n295), .Y(n290) );
  XNOR2XL U227 ( .A(DO_DAC0[2]), .B(DAC1_V[1]), .Y(n292) );
  XNOR2XL U228 ( .A(n307), .B(n308), .Y(N572) );
  XNOR2XL U229 ( .A(n309), .B(n310), .Y(n308) );
  XNOR2XL U230 ( .A(n312), .B(n313), .Y(n307) );
  XNOR2XL U231 ( .A(DAC1_V[8]), .B(TX_EN), .Y(n309) );
  OAI2B11X1 U232 ( .D(sram_rdat[1]), .C(n207), .A(n208), .B(n217), .Y(
        memdatai[1]) );
  AOI22X1 U233 ( .A(regx_rdat[1]), .B(n210), .C(ictlr_inst[1]), .D(n5), .Y(
        n217) );
  OAI211X1 U234 ( .C(n159), .D(n207), .A(n208), .B(n214), .Y(memdatai[4]) );
  AOI22X1 U235 ( .A(regx_rdat[4]), .B(n210), .C(ictlr_inst[4]), .D(n5), .Y(
        n214) );
  OAI211X1 U236 ( .C(n158), .D(n207), .A(n208), .B(n213), .Y(memdatai[5]) );
  AOI22X1 U237 ( .A(regx_rdat[5]), .B(n210), .C(ictlr_inst[5]), .D(n5), .Y(
        n213) );
  OAI211X1 U238 ( .C(n157), .D(n207), .A(n208), .B(n212), .Y(memdatai[6]) );
  AOI22X1 U239 ( .A(regx_rdat[6]), .B(n210), .C(ictlr_inst[6]), .D(n6), .Y(
        n212) );
  OAI211X1 U240 ( .C(n160), .D(n207), .A(n208), .B(n215), .Y(memdatai[3]) );
  AOI22X1 U241 ( .A(regx_rdat[3]), .B(n210), .C(ictlr_inst[3]), .D(n5), .Y(
        n215) );
  OAI211X1 U242 ( .C(n161), .D(n207), .A(n208), .B(n216), .Y(memdatai[2]) );
  AOI22X1 U243 ( .A(regx_rdat[2]), .B(n210), .C(ictlr_inst[2]), .D(n6), .Y(
        n216) );
  OAI2B11X1 U244 ( .D(sram_rdat[0]), .C(n207), .A(n208), .B(n218), .Y(
        memdatai[0]) );
  AOI22X1 U245 ( .A(regx_rdat[0]), .B(n210), .C(ictlr_inst[0]), .D(n6), .Y(
        n218) );
  AO22X1 U246 ( .A(xram_a[8]), .B(n4), .C(iram_a[8]), .D(n10), .Y(SRAM_A[8])
         );
  AO22XL U247 ( .A(xram_a[1]), .B(xram_ce), .C(iram_a[1]), .D(iram_ce), .Y(
        SRAM_A[1]) );
  AO22X1 U248 ( .A(xram_a[10]), .B(n4), .C(iram_a[10]), .D(n10), .Y(SRAM_A[10]) );
  XNOR2XL U249 ( .A(n331), .B(n332), .Y(N1493) );
  XNOR2XL U250 ( .A(DAC1_V[3]), .B(n333), .Y(n332) );
  XNOR2XL U251 ( .A(n334), .B(SRAM_A[9]), .Y(n331) );
  XNOR2XL U252 ( .A(DO_DAC0[4]), .B(n529), .Y(n333) );
  XNOR2XL U253 ( .A(n256), .B(n257), .Y(N586) );
  XNOR2XL U254 ( .A(n258), .B(n259), .Y(n257) );
  XNOR2XL U255 ( .A(n260), .B(SRAM_A[0]), .Y(n256) );
  XNOR2XL U256 ( .A(DO_PWR_I[0]), .B(DO_GPIO[0]), .Y(n258) );
  XNOR2XL U257 ( .A(n261), .B(n262), .Y(N585) );
  XNOR2XL U258 ( .A(n263), .B(n264), .Y(n262) );
  XNOR2XL U259 ( .A(n265), .B(SRAM_A[1]), .Y(n261) );
  XNOR2XL U260 ( .A(DO_PWR_I[1]), .B(DO_GPIO[1]), .Y(n263) );
  XNOR2XL U261 ( .A(n339), .B(n340), .Y(N1488) );
  XNOR2XL U262 ( .A(DAC1_V[4]), .B(n341), .Y(n340) );
  XNOR2XL U263 ( .A(n342), .B(SRAM_A[10]), .Y(n339) );
  XNOR2XL U264 ( .A(DO_DAC0[5]), .B(n530), .Y(n341) );
  XNOR2XL U265 ( .A(n322), .B(n323), .Y(N1498) );
  XNOR2XL U266 ( .A(DAC1_V[2]), .B(n324), .Y(n323) );
  XNOR2XL U267 ( .A(n325), .B(SRAM_A[8]), .Y(n322) );
  XNOR2XL U268 ( .A(DO_DAC0[3]), .B(n528), .Y(n324) );
  XOR2X1 U269 ( .A(n253), .B(SRAM_D[6]), .Y(n342) );
  XNOR2XL U270 ( .A(n347), .B(n348), .Y(N1483) );
  XNOR2XL U271 ( .A(DO_DAC0[6]), .B(n349), .Y(n348) );
  XNOR2XL U272 ( .A(n350), .B(SRAM_D[7]), .Y(n347) );
  XNOR2XL U273 ( .A(n139), .B(dacmux_sel[11]), .Y(n349) );
  ENOX1 U274 ( .A(n127), .B(n119), .C(iram_d[6]), .D(iram_we), .Y(SRAM_D[6])
         );
  ENOX1 U275 ( .A(n128), .B(n119), .C(iram_we), .D(iram_d[7]), .Y(SRAM_D[7])
         );
  XNOR2XL U276 ( .A(n242), .B(n254), .Y(n334) );
  OAI22X1 U277 ( .A(n167), .B(n125), .C(n43), .D(n118), .Y(r_cvcwdat[4]) );
  INVX1 U278 ( .A(xram_d[4]), .Y(n125) );
  OAI22X1 U279 ( .A(n167), .B(n126), .C(n46), .D(n118), .Y(r_cvcwdat[5]) );
  INVX1 U280 ( .A(xram_d[5]), .Y(n126) );
  OAI22AX1 U281 ( .D(xram_d[0]), .C(n167), .A(n118), .B(n33), .Y(r_cvcwdat[0])
         );
  AOI22XL U282 ( .A(xram_d[5]), .B(xram_we), .C(iram_d[5]), .D(iram_we), .Y(
        n242) );
  XNOR2XL U283 ( .A(n243), .B(n255), .Y(n325) );
  ENOXL U284 ( .A(n123), .B(n119), .C(iram_d[3]), .D(iram_we), .Y(SRAM_D[3])
         );
  AOI22X1 U285 ( .A(xram_d[4]), .B(xram_we), .C(iram_d[4]), .D(iram_we), .Y(
        n243) );
  ENOX1 U286 ( .A(n121), .B(n119), .C(iram_d[2]), .D(iram_we), .Y(SRAM_D[2])
         );
  AOI22X1 U287 ( .A(xram_d[0]), .B(xram_we), .C(iram_d[0]), .D(iram_we), .Y(
        n244) );
  ENOX1 U288 ( .A(n120), .B(n119), .C(iram_d[1]), .D(iram_we), .Y(SRAM_D[1])
         );
  NOR21XL U289 ( .B(hit_xr), .A(n5), .Y(n210) );
  INVX1 U290 ( .A(n158), .Y(n140) );
  INVX1 U291 ( .A(n159), .Y(n142) );
  INVX1 U292 ( .A(n157), .Y(n138) );
  INVX1 U293 ( .A(n156), .Y(n136) );
  INVX1 U294 ( .A(n160), .Y(n145) );
  INVX1 U295 ( .A(n161), .Y(n147) );
  OR2X1 U296 ( .A(hit_xr), .B(n6), .Y(n207) );
  XNOR2XL U297 ( .A(n296), .B(n297), .Y(N574) );
  XNOR2XL U298 ( .A(DO_DAC0[7]), .B(n298), .Y(n297) );
  XNOR2XL U299 ( .A(n130), .B(n299), .Y(n296) );
  XNOR2XL U300 ( .A(r_xana_19), .B(n531), .Y(n298) );
  AOI221XL U301 ( .A(n402), .B(pwm_o[0]), .C(n515), .D(r_osc_stop), .E(n423), 
        .Y(n422) );
  OAI22X1 U302 ( .A(n573), .B(n516), .C(n411), .D(n554), .Y(n423) );
  INVX1 U303 ( .A(xram_d[1]), .Y(n120) );
  INVX1 U304 ( .A(xram_d[7]), .Y(n128) );
  INVX1 U305 ( .A(xram_d[6]), .Y(n127) );
  INVX1 U306 ( .A(xram_d[2]), .Y(n121) );
  INVX1 U307 ( .A(xram_d[3]), .Y(n123) );
  XNOR2XL U308 ( .A(DO_DAC0[8]), .B(n532), .Y(n303) );
  XNOR2XL U309 ( .A(dacmux_sel[6]), .B(DO_PWR_I[6]), .Y(n288) );
  XNOR2XL U310 ( .A(dacmux_sel[5]), .B(DO_PWR_I[5]), .Y(n283) );
  XNOR2XL U311 ( .A(dacmux_sel[7]), .B(DO_PWR_I[7]), .Y(n293) );
  XNOR2XL U312 ( .A(o_dodat0_15_), .B(dacmux_sel[15]), .Y(n317) );
  XNOR2XL U313 ( .A(dacmux_sel[16]), .B(dacmux_sel[0]), .Y(n259) );
  XNOR2XL U314 ( .A(dacmux_sel[1]), .B(dacmux_sel[17]), .Y(n264) );
  XNOR2XL U315 ( .A(dacmux_sel[14]), .B(DO_DAC0[9]), .Y(n310) );
  XNOR2XL U316 ( .A(n301), .B(n302), .Y(N573) );
  XNOR2XL U317 ( .A(n304), .B(n305), .Y(n301) );
  XNOR2XL U318 ( .A(DAC1_V[7]), .B(n303), .Y(n302) );
  XNOR2XL U319 ( .A(n306), .B(n250), .Y(n304) );
  XNOR2XL U320 ( .A(n314), .B(n315), .Y(N571) );
  XNOR2XL U321 ( .A(n318), .B(n319), .Y(n314) );
  XNOR2XL U322 ( .A(n316), .B(n317), .Y(n315) );
  XNOR2XL U323 ( .A(n320), .B(n321), .Y(n318) );
  INVX1 U324 ( .A(n168), .Y(n593) );
  NOR2X1 U325 ( .A(n533), .B(n525), .Y(N570) );
  INVX1 U326 ( .A(n172), .Y(n598) );
  INVX1 U327 ( .A(n171), .Y(n592) );
  INVX1 U328 ( .A(n173), .Y(n599) );
  INVX1 U329 ( .A(n170), .Y(n600) );
  INVX1 U330 ( .A(n169), .Y(n597) );
  INVX1 U331 ( .A(pwm_o[0]), .Y(n135) );
  OAI22X1 U332 ( .A(n162), .B(n357), .C(mcuo_scl), .D(n151), .Y(n338) );
  NOR2X1 U333 ( .A(n611), .B(n608), .Y(N610) );
  NOR2X1 U334 ( .A(n621), .B(n618), .Y(N644) );
  NOR2X1 U335 ( .A(n614), .B(n613), .Y(N603) );
  NOR2X1 U336 ( .A(n624), .B(n623), .Y(N637) );
  NOR2X1 U337 ( .A(n615), .B(n614), .Y(N604) );
  NOR2X1 U338 ( .A(n625), .B(n624), .Y(N638) );
  NOR2X1 U339 ( .A(n611), .B(n609), .Y(N598) );
  NOR2X1 U340 ( .A(n621), .B(n619), .Y(N632) );
  NOR2X1 U341 ( .A(n610), .B(n609), .Y(N597) );
  NOR2X1 U342 ( .A(n620), .B(n619), .Y(N631) );
  NOR2X1 U343 ( .A(n615), .B(n608), .Y(N608) );
  NOR2X1 U344 ( .A(n625), .B(n618), .Y(N642) );
  INVX1 U345 ( .A(n177), .Y(n588) );
  AOI221XL U346 ( .A(N635), .B(n13), .C(N601), .D(n569), .E(n597), .Y(n453) );
  NOR2X1 U347 ( .A(n612), .B(n610), .Y(N601) );
  NOR2X1 U348 ( .A(n622), .B(n620), .Y(N635) );
  AOI221XL U349 ( .A(N639), .B(n13), .C(N605), .D(n569), .E(n591), .Y(n470) );
  NOR2X1 U350 ( .A(n614), .B(n610), .Y(N605) );
  NOR2X1 U351 ( .A(n624), .B(n620), .Y(N639) );
  AOI221XL U352 ( .A(N636), .B(n13), .C(N602), .D(n569), .E(n593), .Y(n459) );
  NOR2X1 U353 ( .A(n612), .B(n611), .Y(N602) );
  NOR2X1 U354 ( .A(n622), .B(n621), .Y(N636) );
  NAND2X1 U355 ( .A(n472), .B(n470), .Y(n448) );
  NOR2X1 U356 ( .A(n615), .B(n612), .Y(N600) );
  NOR2X1 U357 ( .A(n625), .B(n622), .Y(N634) );
  NOR2X1 U358 ( .A(n613), .B(n609), .Y(N596) );
  NOR2X1 U359 ( .A(n623), .B(n619), .Y(N629) );
  NOR2X1 U360 ( .A(n613), .B(n612), .Y(N599) );
  NOR2X1 U361 ( .A(n623), .B(n622), .Y(N633) );
  NOR2X1 U362 ( .A(n613), .B(n608), .Y(N607) );
  NOR2X1 U363 ( .A(n623), .B(n618), .Y(N641) );
  NOR2X1 U364 ( .A(n614), .B(n611), .Y(N606) );
  NOR2X1 U365 ( .A(n624), .B(n621), .Y(N640) );
  INVX1 U366 ( .A(n240), .Y(n134) );
  INVX1 U367 ( .A(n330), .Y(do_opt_1) );
  NOR2X1 U368 ( .A(n70), .B(n254), .Y(OE_GPIO[1]) );
  NOR2X1 U369 ( .A(n71), .B(n255), .Y(OE_GPIO[0]) );
  NOR2X1 U370 ( .A(n70), .B(n251), .Y(OE_GPIO[4]) );
  NOR2X1 U371 ( .A(n71), .B(n252), .Y(OE_GPIO[3]) );
  NOR2X1 U372 ( .A(n70), .B(n253), .Y(OE_GPIO[2]) );
  NAND2X1 U373 ( .A(n249), .B(n74), .Y(OE_GPIO[6]) );
  NAND2X1 U374 ( .A(n250), .B(n78), .Y(OE_GPIO[5]) );
  INVX1 U375 ( .A(n181), .Y(n596) );
  INVX1 U376 ( .A(n182), .Y(n590) );
  INVX1 U377 ( .A(n189), .Y(n151) );
  INVX1 U378 ( .A(n176), .Y(n595) );
  INVX1 U379 ( .A(n180), .Y(n591) );
  AO222X1 U380 ( .A(di_xanav[1]), .B(n436), .C(di_xanav[0]), .D(n440), .E(n580), .F(n435), .Y(n442) );
  NAND31X1 U381 ( .C(n488), .A(n472), .B(n453), .Y(n496) );
  XNOR2XL U382 ( .A(DAC3_V[1]), .B(n522), .Y(n265) );
  AOI222XL U383 ( .A(n188), .B(n196), .C(n197), .D(n189), .E(n150), .F(n198), 
        .Y(n507) );
  INVX1 U384 ( .A(n393), .Y(n586) );
  OAI22X1 U385 ( .A(n443), .B(n453), .C(n454), .D(n455), .Y(n452) );
  OAI21X1 U386 ( .B(do_opt_1), .C(n549), .A(n548), .Y(n345) );
  NOR3XL U387 ( .A(n188), .B(n183), .C(n451), .Y(di_cc) );
  INVX1 U388 ( .A(n418), .Y(n581) );
  AOI21X1 U389 ( .B(n455), .C(n456), .A(n451), .Y(n479) );
  INVX1 U390 ( .A(n443), .Y(n580) );
  INVX1 U391 ( .A(n472), .Y(n562) );
  AOI222XL U392 ( .A(n188), .B(n184), .C(n189), .D(n186), .E(n150), .F(n187), 
        .Y(n505) );
  INVX1 U393 ( .A(n179), .Y(n589) );
  INVX1 U394 ( .A(n178), .Y(n594) );
  INVX1 U395 ( .A(n185), .Y(n162) );
  INVX1 U396 ( .A(n451), .Y(n584) );
  AOI222XL U397 ( .A(n183), .B(n196), .C(n197), .D(n185), .E(n155), .F(n198), 
        .Y(n506) );
  AOI222XL U398 ( .A(n183), .B(n184), .C(n185), .D(n186), .E(n155), .F(n187), 
        .Y(n504) );
  INVX1 U399 ( .A(n321), .Y(TX_DAT) );
  INVX1 U400 ( .A(n388), .Y(n582) );
  INVX1 U401 ( .A(n389), .Y(n583) );
  INVX1 U402 ( .A(di_gpio[0]), .Y(n133) );
  INVX1 U403 ( .A(n311), .Y(n534) );
  INVX1 U404 ( .A(n438), .Y(n143) );
  INVX1 U405 ( .A(n440), .Y(n144) );
  INVX1 U406 ( .A(n437), .Y(n585) );
  INVX1 U407 ( .A(n454), .Y(n587) );
  XNOR2XL U408 ( .A(DO_DAC0[10]), .B(DAC1_V[9]), .Y(n316) );
  XOR2X1 U409 ( .A(DAC1_V[5]), .B(n252), .Y(n350) );
  XNOR2XL U410 ( .A(DAC1_V[6]), .B(n251), .Y(n299) );
  OAI22X1 U411 ( .A(n129), .B(n380), .C(n135), .D(n381), .Y(n379) );
  AOI221XL U412 ( .A(n402), .B(pwm_o[1]), .C(n515), .D(o_dodat0_15_), .E(n410), 
        .Y(n409) );
  OAI22X1 U413 ( .A(n516), .B(n544), .C(n555), .D(n411), .Y(n410) );
  OAI22X1 U414 ( .A(n153), .B(n357), .C(mcuo_scl), .D(n149), .Y(n501) );
  AOI221XL U415 ( .A(n519), .B(CC1_DOB), .C(n412), .D(n523), .E(n424), .Y(n421) );
  OAI32X1 U416 ( .A(n518), .B(n521), .C(n555), .D(n414), .E(n131), .Y(n424) );
  AOI221XL U417 ( .A(n519), .B(CC2_DOB), .C(n412), .D(n522), .E(n413), .Y(n408) );
  OAI22X1 U418 ( .A(n414), .B(n141), .C(n520), .D(n518), .Y(n413) );
  INVX1 U419 ( .A(n279), .Y(CC2_DOB) );
  AND2X1 U420 ( .A(n77), .B(n109), .Y(i2c_ev_6_) );
  INVX1 U421 ( .A(r_ocdrv_enz), .Y(n554) );
  OAI22X1 U422 ( .A(n396), .B(n357), .C(mcuo_scl), .D(n397), .Y(n362) );
  INVX1 U423 ( .A(n183), .Y(n153) );
  INVX1 U424 ( .A(n188), .Y(n149) );
  NAND2X1 U425 ( .A(n542), .B(n508), .Y(n381) );
  AOI221XL U426 ( .A(n519), .B(di_pro[5]), .C(n412), .D(n587), .E(n417), .Y(
        n415) );
  OAI22X1 U427 ( .A(n418), .B(n414), .C(n389), .D(n518), .Y(n417) );
  INVX1 U428 ( .A(n425), .Y(n523) );
  INVX1 U429 ( .A(n375), .Y(n522) );
  INVX1 U430 ( .A(n411), .Y(n519) );
  INVX1 U431 ( .A(n402), .Y(n518) );
  INVX1 U432 ( .A(n376), .Y(n211) );
  INVX1 U433 ( .A(n414), .Y(n515) );
  INVX1 U434 ( .A(n374), .Y(n512) );
  INVX1 U435 ( .A(n412), .Y(n516) );
  NOR2X1 U436 ( .A(n311), .B(n69), .Y(TX_EN) );
  INVX1 U437 ( .A(n380), .Y(n511) );
  INVX1 U438 ( .A(n397), .Y(n150) );
  INVX1 U439 ( .A(n396), .Y(n155) );
  INVX1 U440 ( .A(o_dodat5_2_), .Y(n137) );
  INVX1 U441 ( .A(sh_hold), .Y(n525) );
  INVX1 U442 ( .A(n430), .Y(n124) );
  INVX1 U443 ( .A(n241), .Y(n122) );
  NOR21XL U444 ( .B(dacmux_sel[5]), .A(n55), .Y(SAMPL_SEL[5]) );
  NOR21XL U445 ( .B(dacmux_sel[4]), .A(n55), .Y(SAMPL_SEL[4]) );
  NOR21XL U446 ( .B(dacmux_sel[6]), .A(n55), .Y(SAMPL_SEL[6]) );
  NOR21XL U447 ( .B(dacmux_sel[7]), .A(n55), .Y(SAMPL_SEL[7]) );
  NOR21XL U448 ( .B(dacmux_sel[1]), .A(n55), .Y(SAMPL_SEL[1]) );
  NOR21XL U449 ( .B(dacmux_sel[14]), .A(n56), .Y(SAMPL_SEL[14]) );
  NOR21XL U450 ( .B(dacmux_sel[15]), .A(n56), .Y(SAMPL_SEL[15]) );
  NOR21XL U451 ( .B(dacmux_sel[16]), .A(n56), .Y(SAMPL_SEL[16]) );
  NOR21XL U452 ( .B(dacmux_sel[17]), .A(n55), .Y(SAMPL_SEL[17]) );
  NOR21XL U453 ( .B(dacmux_sel[0]), .A(n56), .Y(SAMPL_SEL[0]) );
  NOR21XL U454 ( .B(r_xana_19), .A(n55), .Y(STB_RP) );
  NOR21XL U455 ( .B(n305), .A(n67), .Y(DO_VOOC[1]) );
  NOR21XL U456 ( .B(n313), .A(n67), .Y(DO_VOOC[2]) );
  NOR21XL U457 ( .B(n320), .A(n66), .Y(DO_VOOC[3]) );
  NOR21XL U458 ( .B(PWRDN), .A(n521), .Y(VPP_0V) );
  OR2X2 U459 ( .A(pmem_csb), .B(n73), .Y(PMEM_CSB) );
  NAND2X1 U460 ( .A(N630), .B(n499), .Y(n154) );
  NOR2X1 U461 ( .A(n625), .B(n619), .Y(N630) );
  NAND2X1 U462 ( .A(sll_223_2_A_0_), .B(n604), .Y(N595) );
  NAND2X1 U463 ( .A(n603), .B(n577), .Y(n619) );
  NAND2X1 U464 ( .A(n601), .B(n616), .Y(n620) );
  NAND2X1 U465 ( .A(n579), .B(n606), .Y(n610) );
  NAND2X1 U466 ( .A(n602), .B(n617), .Y(n625) );
  NOR2X1 U467 ( .A(n70), .B(n575), .Y(PMEM_CLK[0]) );
  NOR2X1 U468 ( .A(n69), .B(n574), .Y(PMEM_CLK[1]) );
  NAND3X1 U469 ( .A(n606), .B(n607), .C(N595), .Y(n613) );
  NAND3X1 U470 ( .A(n616), .B(n617), .C(sll_223_2_A_0_), .Y(n623) );
  AND2X1 U471 ( .A(dacmux_sel[11]), .B(n93), .Y(SAMPL_SEL[11]) );
  NAND2X1 U472 ( .A(n603), .B(n577), .Y(n609) );
  NAND2X1 U473 ( .A(n578), .B(n607), .Y(n615) );
  INVX1 U474 ( .A(atpg_en), .Y(n92) );
  INVX1 U475 ( .A(atpg_en), .Y(n93) );
  INVX1 U476 ( .A(atpg_en), .Y(n94) );
  NOR2X1 U477 ( .A(n555), .B(n69), .Y(PWRDN) );
  NOR2X1 U478 ( .A(n72), .B(n604), .Y(lt_gpi[0]) );
  NOR2X1 U479 ( .A(n69), .B(n375), .Y(DO_SRCCTL[4]) );
  NOR2X1 U480 ( .A(n69), .B(n425), .Y(DO_SRCCTL[1]) );
  NOR2X1 U481 ( .A(n71), .B(n141), .Y(ANA_REGX[12]) );
  NOR2X1 U482 ( .A(n71), .B(n533), .Y(SH_RST) );
  NOR2X1 U483 ( .A(n70), .B(n130), .Y(DO_VOOC[0]) );
  NOR2X1 U484 ( .A(n71), .B(n520), .Y(VPP_SEL) );
  NOR2X1 U485 ( .A(n69), .B(n131), .Y(DO_SRCCTL[0]) );
  NOR2X1 U486 ( .A(n71), .B(n529), .Y(SAMPL_SEL[9]) );
  NOR2X1 U487 ( .A(n71), .B(n528), .Y(SAMPL_SEL[8]) );
  NOR2X1 U488 ( .A(n70), .B(n531), .Y(SAMPL_SEL[12]) );
  NOR2X1 U489 ( .A(n71), .B(n526), .Y(SAMPL_SEL[2]) );
  NOR2X1 U490 ( .A(n71), .B(n527), .Y(SAMPL_SEL[3]) );
  NOR2X1 U491 ( .A(n70), .B(n532), .Y(SAMPL_SEL[13]) );
  NOR2X1 U492 ( .A(n70), .B(n530), .Y(SAMPL_SEL[10]) );
  NOR2X1 U493 ( .A(n69), .B(n539), .Y(DO_SRCCTL[5]) );
  NOR2X1 U494 ( .A(n69), .B(n541), .Y(DO_DPDN[3]) );
  NOR2X1 U495 ( .A(n70), .B(n536), .Y(DO_CCCTL[0]) );
  NOR2X1 U496 ( .A(n72), .B(n306), .Y(ANAOPT[5]) );
  INVX1 U497 ( .A(n616), .Y(n602) );
  INVX1 U498 ( .A(n606), .Y(n578) );
  INVX1 U499 ( .A(n617), .Y(n601) );
  INVX1 U500 ( .A(n607), .Y(n579) );
  NAND2X1 U501 ( .A(n139), .B(n76), .Y(RD_ENB) );
  NAND2X1 U502 ( .A(n544), .B(n75), .Y(SLEEP) );
  OAI22AX1 U503 ( .D(r_do_ts[6]), .C(n431), .A(r_do_ts[6]), .B(n432), .Y(n295)
         );
  EORX1 U504 ( .A(r_do_ts[3]), .B(n433), .C(r_do_ts[3]), .D(n434), .Y(n432) );
  AOI22AXL U505 ( .A(r_do_ts[3]), .B(n441), .D(r_do_ts[3]), .C(n442), .Y(n431)
         );
  OAI211X1 U506 ( .C(n437), .D(n438), .A(n144), .B(n439), .Y(n433) );
  NAND4X1 U507 ( .A(n474), .B(n475), .C(n476), .D(n477), .Y(DO_GPIO[4]) );
  AOI221XL U508 ( .A(n464), .B(n583), .C(mcu_dbgpo[18]), .D(n478), .E(n479), 
        .Y(n477) );
  AOI222XL U509 ( .A(upd_dbgpo[18]), .B(n558), .C(n449), .D(n480), .E(n563), 
        .F(n534), .Y(n476) );
  AOI222XL U510 ( .A(comp_smpl[1]), .B(n568), .C(slvo_sda), .D(n567), .E(
        r_dpdmctl[4]), .F(n564), .Y(n475) );
  INVX1 U511 ( .A(pmem_clk[1]), .Y(n574) );
  AO22X1 U512 ( .A(xram_a[7]), .B(xram_ce), .C(iram_a[7]), .D(iram_ce), .Y(
        SRAM_A[7]) );
  AO22X1 U513 ( .A(n4), .B(xram_a[9]), .C(n10), .D(iram_a[9]), .Y(SRAM_A[9])
         );
  OR2X1 U514 ( .A(slvo_early), .B(slvo_re), .Y(n77) );
  NOR21XL U515 ( .B(n109), .A(n108), .Y(sse_prefetch) );
  AND4X1 U516 ( .A(r_pg0_sel[2]), .B(r_pg0_sel[3]), .C(n107), .D(n106), .Y(
        n108) );
  INVX1 U517 ( .A(r_pg0_sel[1]), .Y(n106) );
  INVX1 U518 ( .A(r_pg0_sel[0]), .Y(n107) );
  INVX1 U519 ( .A(sse_adr[7]), .Y(n109) );
  AOI221XL U520 ( .A(r_accctl[4]), .B(n564), .C(comp_smpl[3]), .D(n568), .E(
        n457), .Y(n445) );
  OAI22X1 U521 ( .A(n458), .B(n536), .C(n418), .D(n459), .Y(n457) );
  OAI31XL U522 ( .A(n205), .B(o_cpurst), .C(hit_ps), .D(n206), .Y(mempsack) );
  NOR2X1 U523 ( .A(mempsrd), .B(mempswr), .Y(n205) );
  NAND2X1 U524 ( .A(ictlr_psack), .B(hit_ps), .Y(n206) );
  AOI22X1 U525 ( .A(comp_smpl[0]), .B(n568), .C(r_vpp_en), .D(n560), .Y(n483)
         );
  NAND4X1 U526 ( .A(n483), .B(n484), .C(n485), .D(n486), .Y(DO_GPIO[3]) );
  AOI22X1 U527 ( .A(n567), .B(n585), .C(n556), .D(n584), .Y(n484) );
  AOI222XL U528 ( .A(mcu_dbgpo[16]), .B(n448), .C(n464), .D(di_pro[0]), .E(
        prx_rcvinf[4]), .F(n465), .Y(n486) );
  AOI22X1 U529 ( .A(N449), .B(n487), .C(mcu_dbgpo[21]), .D(n488), .Y(n485) );
  NAND4X1 U530 ( .A(n460), .B(n461), .C(n462), .D(n463), .Y(DO_GPIO[5]) );
  AOI222XL U531 ( .A(n563), .B(TX_DAT), .C(n576), .D(i_rstz), .E(n556), .F(
        dp_comp), .Y(n462) );
  AOI222XL U532 ( .A(mcu_dbgpo[22]), .B(n566), .C(fcp_do), .D(n565), .E(
        mcu_dbgpo[19]), .F(n562), .Y(n460) );
  AOI221XL U533 ( .A(n464), .B(n582), .C(upd_dbgpo[17]), .D(n465), .E(n466), 
        .Y(n463) );
  NAND4X1 U534 ( .A(n444), .B(n445), .C(n446), .D(n447), .Y(DO_GPIO[6]) );
  AOI221XL U535 ( .A(n559), .B(n584), .C(n567), .D(TX_DAT), .E(n452), .Y(n446)
         );
  AOI222XL U536 ( .A(mcu_dbgpo[16]), .B(n566), .C(pmem_pgm), .D(n560), .E(
        fcp_oe), .F(n565), .Y(n444) );
  AOI221XL U537 ( .A(mcu_dbgpo[17]), .B(n448), .C(do_p0[6]), .D(n449), .E(n450), .Y(n447) );
  AOI221XL U538 ( .A(comp_smpl[2]), .B(n568), .C(pmem_re), .D(n560), .E(n469), 
        .Y(n461) );
  OAI22X1 U539 ( .A(n470), .B(n129), .C(n471), .D(n541), .Y(n469) );
  AOI21X1 U540 ( .B(SRAM_RDAT[7]), .C(n87), .A(n593), .Y(n156) );
  OAI21BBX1 U541 ( .A(SRAM_RDAT[0]), .B(n81), .C(n175), .Y(sram_rdat[0]) );
  OAI21BBX1 U542 ( .A(SRAM_RDAT[1]), .B(n80), .C(n174), .Y(sram_rdat[1]) );
  AOI21X1 U543 ( .B(SRAM_RDAT[5]), .C(n87), .A(n600), .Y(n158) );
  AOI21X1 U544 ( .B(SRAM_RDAT[6]), .C(n88), .A(n597), .Y(n157) );
  AOI21X1 U545 ( .B(SRAM_RDAT[4]), .C(n88), .A(n592), .Y(n159) );
  AOI21X1 U546 ( .B(SRAM_RDAT[3]), .C(n86), .A(n598), .Y(n160) );
  AOI21X1 U547 ( .B(SRAM_RDAT[2]), .C(n87), .A(n599), .Y(n161) );
  OAI21BBX1 U548 ( .A(hit_ps), .B(mempsrd), .C(n5), .Y(n208) );
  INVX1 U549 ( .A(n398), .Y(n130) );
  OAI221X1 U550 ( .A(r_dpdmctl[0]), .B(n399), .C(n400), .D(n543), .E(n401), 
        .Y(n398) );
  INVX1 U551 ( .A(r_dpdmctl[0]), .Y(n543) );
  NAND4X1 U552 ( .A(n402), .B(n403), .C(n514), .D(n513), .Y(n401) );
  AOI22X1 U553 ( .A(n419), .B(n513), .C(r_dndo_sel[3]), .D(n420), .Y(n399) );
  OAI21BX1 U554 ( .C(r_dndo_sel[0]), .B(n426), .A(n427), .Y(n419) );
  OAI22X1 U555 ( .A(n421), .B(n514), .C(r_dndo_sel[2]), .D(n422), .Y(n420) );
  AOI33X1 U556 ( .A(n402), .B(di_pro[0]), .C(r_dndo_sel[2]), .D(n534), .E(n514), .F(n412), .Y(n427) );
  INVX1 U557 ( .A(r_osc_gate), .Y(n573) );
  NOR21XL U558 ( .B(esfrm_rrdy), .A(prl_cany0), .Y(sse_rdrdy) );
  NOR21XL U559 ( .B(bist_r_ctl[5]), .A(n55), .Y(SRAM_OEB) );
  INVX1 U560 ( .A(dacmux_sel[12]), .Y(n531) );
  INVX1 U561 ( .A(dacmux_sel[2]), .Y(n526) );
  INVX1 U562 ( .A(dacmux_sel[3]), .Y(n527) );
  INVX1 U563 ( .A(dacmux_sel[13]), .Y(n532) );
  INVX1 U564 ( .A(dacmux_sel[10]), .Y(n530) );
  INVX1 U565 ( .A(dacmux_sel[8]), .Y(n528) );
  INVX1 U566 ( .A(dacmux_sel[9]), .Y(n529) );
  NAND2X1 U567 ( .A(d_dodat[7]), .B(n68), .Y(n168) );
  NAND2X1 U568 ( .A(d_dodat[4]), .B(n67), .Y(n171) );
  NAND2X1 U569 ( .A(d_dodat[2]), .B(n68), .Y(n173) );
  NAND2X1 U570 ( .A(d_dodat[3]), .B(n68), .Y(n172) );
  NAND2X1 U571 ( .A(d_dodat[5]), .B(n68), .Y(n170) );
  NAND2X1 U572 ( .A(d_dodat[6]), .B(n68), .Y(n169) );
  NAND2X1 U573 ( .A(d_dodat[0]), .B(n69), .Y(n175) );
  NAND2X1 U574 ( .A(d_dodat[1]), .B(n68), .Y(n174) );
  INVX1 U575 ( .A(sh_rst), .Y(n533) );
  AND2X1 U576 ( .A(esfrm_rrdy), .B(prl_cany0), .Y(upd_rdrdy) );
  XNOR2XL U577 ( .A(do_p0[4]), .B(n135), .Y(n480) );
  OAI22X1 U578 ( .A(n311), .B(n467), .C(n468), .D(n557), .Y(n466) );
  XNOR2XL U579 ( .A(pwm_o[1]), .B(do_p0[5]), .Y(n468) );
  NOR2X1 U580 ( .A(n610), .B(n608), .Y(N609) );
  NOR2X1 U581 ( .A(n620), .B(n618), .Y(N643) );
  MUX2X1 U582 ( .D0(n111), .D1(n110), .S(N260), .Y(N449) );
  MUX4X1 U583 ( .D0(do_p0[2]), .D1(do_p0[3]), .D2(do_opt[6]), .D3(do_opt[7]), 
        .S0(N258), .S1(N259), .Y(n110) );
  MUX4X1 U584 ( .D0(do_opt_0), .D1(do_opt_1), .D2(do_p0[0]), .D3(do_p0[1]), 
        .S0(N258), .S1(N259), .Y(n111) );
  MUX2X1 U585 ( .D0(n113), .D1(n112), .S(N263), .Y(N450) );
  MUX4X1 U586 ( .D0(do_p0[2]), .D1(do_p0[3]), .D2(do_opt[6]), .D3(do_opt[7]), 
        .S0(N261), .S1(N262), .Y(n112) );
  MUX4X1 U587 ( .D0(do_opt_0), .D1(do_opt_1), .D2(do_p0[0]), .D3(do_p0[1]), 
        .S0(N261), .S1(N262), .Y(n113) );
  OR2X1 U588 ( .A(mcu_ram_r), .B(mcu_ram_w), .Y(ramacc) );
  INVX1 U589 ( .A(n500), .Y(n569) );
  OAI211X1 U590 ( .C(di_tst), .D(r_gpio_tm), .A(i_rstz), .B(n86), .Y(n500) );
  OAI21X1 U591 ( .B(hwi2c_stretch), .C(pmem_pgm), .A(r_strtch), .Y(n357) );
  OAI22X1 U592 ( .A(slvo_sda), .B(n162), .C(mcuo_sda), .D(n151), .Y(n330) );
  AOI21X1 U593 ( .B(DI_GPIO[3]), .C(n87), .A(n598), .Y(n240) );
  MUX2X1 U594 ( .D0(n117), .D1(n116), .S(N269), .Y(DO_GPIO[0]) );
  MUX4X1 U595 ( .D0(do_p0[2]), .D1(do_p0[3]), .D2(do_opt[6]), .D3(do_opt[7]), 
        .S0(N267), .S1(N268), .Y(n116) );
  MUX4X1 U596 ( .D0(do_opt_0), .D1(do_opt_1), .D2(do_p0[0]), .D3(do_p0[1]), 
        .S0(N267), .S1(N268), .Y(n117) );
  MUX2X1 U597 ( .D0(n115), .D1(n114), .S(N266), .Y(DO_GPIO[1]) );
  MUX4X1 U598 ( .D0(do_p0[2]), .D1(do_p0[3]), .D2(do_opt[6]), .D3(do_opt[7]), 
        .S0(N264), .S1(N265), .Y(n114) );
  MUX4X1 U599 ( .D0(do_opt_0), .D1(do_opt_1), .D2(do_p0[0]), .D3(do_p0[1]), 
        .S0(N264), .S1(N265), .Y(n115) );
  AND3X1 U600 ( .A(n352), .B(i_rstz), .C(n353), .Y(n300) );
  NAND2X1 U601 ( .A(d_dodat[13]), .B(n69), .Y(n177) );
  OAI21X1 U602 ( .B(n343), .C(n300), .A(n327), .Y(n253) );
  NOR21XL U603 ( .B(r_gpio_oe[2]), .A(n344), .Y(n343) );
  AOI221XL U604 ( .A(n338), .B(n549), .C(n345), .D(n547), .E(n346), .Y(n344)
         );
  AOI31X1 U605 ( .A(N261), .B(n570), .C(N262), .D(n547), .Y(n346) );
  OAI21X1 U606 ( .B(n351), .C(n300), .A(n327), .Y(n252) );
  NOR21XL U607 ( .B(r_gpio_oe[3]), .A(n354), .Y(n351) );
  AOI221XL U608 ( .A(n338), .B(n546), .C(n355), .D(n545), .E(n356), .Y(n354)
         );
  AOI31X1 U609 ( .A(N258), .B(n570), .C(N259), .D(n545), .Y(n356) );
  NOR2X1 U610 ( .A(r_i2cmcu_route[0]), .B(r_i2cmcu_route[1]), .Y(n189) );
  NAND2X1 U611 ( .A(d_dodat[15]), .B(n68), .Y(n176) );
  NAND2X1 U612 ( .A(d_dodat[8]), .B(n67), .Y(n182) );
  NAND2X1 U613 ( .A(d_dodat[9]), .B(n68), .Y(n181) );
  NAND2X1 U614 ( .A(d_dodat[10]), .B(n68), .Y(n180) );
  OAI22AX1 U615 ( .D(n220), .C(n221), .A(n133), .B(n220), .Y(exint[1]) );
  NAND3X1 U616 ( .A(N267), .B(n552), .C(N269), .Y(n220) );
  AOI22AXL U617 ( .A(n222), .B(n223), .D(n223), .C(di_gpio[1]), .Y(n221) );
  NAND3X1 U618 ( .A(N264), .B(n550), .C(N266), .Y(n223) );
  NOR3XL U619 ( .A(r_gpio_oe[5]), .B(n561), .C(n300), .Y(n250) );
  NOR3XL U620 ( .A(r_gpio_oe[6]), .B(n561), .C(n300), .Y(n249) );
  NOR2X1 U621 ( .A(r_gpio_oe[4]), .B(n300), .Y(n251) );
  OAI22AX1 U622 ( .D(n226), .C(n227), .A(n133), .B(n226), .Y(exint[0]) );
  NAND3X1 U623 ( .A(n553), .B(n552), .C(N269), .Y(n226) );
  AOI22AXL U624 ( .A(n228), .B(n229), .D(n229), .C(di_gpio[1]), .Y(n227) );
  NAND3X1 U625 ( .A(n551), .B(n550), .C(N266), .Y(n229) );
  ENOX1 U626 ( .A(n224), .B(n225), .C(di_gpio[2]), .D(n224), .Y(n222) );
  NOR3XL U627 ( .A(n549), .B(N262), .C(n547), .Y(n224) );
  NOR4XL U628 ( .A(N259), .B(n134), .C(n546), .D(n545), .Y(n225) );
  NAND3X1 U629 ( .A(n335), .B(n327), .C(r_gpio_oe[1]), .Y(n254) );
  OAI221X1 U630 ( .A(N266), .B(n336), .C(N264), .D(do_opt_0), .E(n337), .Y(
        n335) );
  OAI31XL U631 ( .A(n550), .B(s0_rxdoe), .C(n551), .D(N266), .Y(n337) );
  AOI21X1 U632 ( .B(N264), .C(n330), .A(N265), .Y(n336) );
  NAND3X1 U633 ( .A(n326), .B(n327), .C(r_gpio_oe[0]), .Y(n255) );
  OAI221X1 U634 ( .A(N269), .B(n328), .C(N267), .D(do_opt_0), .E(n329), .Y(
        n326) );
  OAI31XL U635 ( .A(n552), .B(s0_rxdoe), .C(n553), .D(N269), .Y(n329) );
  AOI21X1 U636 ( .B(N267), .C(n330), .A(N268), .Y(n328) );
  ENOX1 U637 ( .A(n230), .B(n231), .C(di_gpio[2]), .D(n230), .Y(n228) );
  NOR3XL U638 ( .A(N261), .B(N262), .C(n547), .Y(n230) );
  NOR4XL U639 ( .A(N259), .B(N258), .C(n134), .D(n545), .Y(n231) );
  AOI21X1 U640 ( .B(CC1_DI), .C(n93), .A(n593), .Y(n393) );
  AOI21X1 U641 ( .B(SRCI[3]), .C(n87), .A(n591), .Y(n418) );
  AOI21X1 U642 ( .B(RX_DAT), .C(n88), .A(n596), .Y(n451) );
  AOI21X1 U643 ( .B(SRCI[4]), .C(n88), .A(n589), .Y(n443) );
  OAI21BBX1 U644 ( .A(DI_GPIO[1]), .B(n83), .C(n174), .Y(di_gpio[1]) );
  OAI21BBX1 U645 ( .A(DI_GPIO[2]), .B(n83), .C(n173), .Y(di_gpio[2]) );
  AO22X1 U646 ( .A(n558), .B(di_cc), .C(x_clk), .D(n576), .Y(n450) );
  NOR2X1 U647 ( .A(ptx_oe), .B(r_fortxen), .Y(n311) );
  OAI21BBX1 U648 ( .A(DM_COMP), .B(n85), .C(n178), .Y(dm_comp) );
  NOR2X1 U649 ( .A(r_i2cslv_route[0]), .B(r_i2cslv_route[1]), .Y(n185) );
  NAND2X1 U650 ( .A(d_dodat[12]), .B(n67), .Y(n178) );
  NAND2X1 U651 ( .A(d_dodat[11]), .B(n68), .Y(n179) );
  EORX1 U652 ( .A(di_gpio[0]), .B(n190), .C(n190), .D(n191), .Y(n186) );
  NOR3XL U653 ( .A(N268), .B(N269), .C(N267), .Y(n190) );
  AOI22AXL U654 ( .A(n192), .B(di_gpio[1]), .D(n192), .C(n193), .Y(n191) );
  NOR3XL U655 ( .A(N265), .B(N266), .C(N264), .Y(n192) );
  AOI222XL U656 ( .A(n435), .B(dp_comp), .C(n143), .D(n586), .E(divff_5), .F(
        n436), .Y(n434) );
  AOI22X1 U657 ( .A(divff_8), .B(n436), .C(n435), .D(dm_comp), .Y(n439) );
  EORX1 U658 ( .A(di_gpio[0]), .B(n199), .C(n199), .D(n200), .Y(n197) );
  NOR3XL U659 ( .A(N268), .B(N269), .C(n553), .Y(n199) );
  AOI22AXL U660 ( .A(n201), .B(di_gpio[1]), .D(n201), .C(n202), .Y(n200) );
  NOR3XL U661 ( .A(N265), .B(N266), .C(n551), .Y(n201) );
  ENOX1 U662 ( .A(n194), .B(n195), .C(di_gpio[2]), .D(n194), .Y(n193) );
  NOR3XL U663 ( .A(N262), .B(N263), .C(N261), .Y(n194) );
  NOR4XL U664 ( .A(N260), .B(N259), .C(N258), .D(n134), .Y(n195) );
  ENOX1 U665 ( .A(n203), .B(n204), .C(di_gpio[2]), .D(n203), .Y(n202) );
  NOR3XL U666 ( .A(N262), .B(N263), .C(n549), .Y(n203) );
  NOR4XL U667 ( .A(N260), .B(N259), .C(n134), .D(n546), .Y(n204) );
  OAI21AX1 U668 ( .B(do_opt_1), .C(n546), .A(N259), .Y(n355) );
  AOI21X1 U669 ( .B(SRCI[2]), .C(n88), .A(n596), .Y(n388) );
  AOI21X1 U670 ( .B(SRCI[1]), .C(n88), .A(n590), .Y(n389) );
  AOI21X1 U671 ( .B(CC2_DI), .C(n87), .A(n595), .Y(n437) );
  AOI21X1 U672 ( .B(DAC1_COMP), .C(n86), .A(n590), .Y(n454) );
  AOI21X1 U673 ( .B(RX_SQL), .C(n80), .A(n589), .Y(n430) );
  NOR21XL U674 ( .B(r_do_ts[5]), .A(r_do_ts[4]), .Y(n435) );
  NOR21XL U675 ( .B(r_do_ts[4]), .A(r_do_ts[5]), .Y(n436) );
  OAI21BBX1 U676 ( .A(DI_GPIO[0]), .B(n84), .C(n175), .Y(di_gpio[0]) );
  OAI21BBX1 U677 ( .A(SRCI[5]), .B(n86), .C(n178), .Y(di_pro[5]) );
  OAI21BBX1 U678 ( .A(DP_COMP), .B(n85), .C(n177), .Y(dp_comp) );
  NOR2X1 U679 ( .A(n152), .B(r_i2cmcu_route[1]), .Y(n188) );
  NOR2X1 U680 ( .A(n163), .B(r_i2cslv_route[1]), .Y(n183) );
  OAI21BBX1 U681 ( .A(SRCI[0]), .B(n85), .C(n168), .Y(di_pro[0]) );
  OAI21BBX1 U682 ( .A(DM_FAULT), .B(n85), .C(n176), .Y(di_aswk[3]) );
  NOR2X1 U683 ( .A(r_do_ts[4]), .B(r_do_ts[5]), .Y(n440) );
  NAND2X1 U684 ( .A(r_do_ts[5]), .B(r_do_ts[4]), .Y(n438) );
  INVX1 U685 ( .A(N258), .Y(n546) );
  INVX1 U686 ( .A(N265), .Y(n550) );
  INVX1 U687 ( .A(N260), .Y(n545) );
  INVX1 U688 ( .A(N261), .Y(n549) );
  INVX1 U689 ( .A(N267), .Y(n553) );
  OAI21BBX1 U690 ( .A(XANAV[1]), .B(n84), .C(n174), .Y(di_xanav[1]) );
  OAI21BBX1 U691 ( .A(XANAV[0]), .B(n84), .C(n175), .Y(di_xanav[0]) );
  INVX1 U692 ( .A(N264), .Y(n551) );
  INVX1 U693 ( .A(N263), .Y(n547) );
  INVX1 U694 ( .A(N268), .Y(n552) );
  INVX1 U695 ( .A(r_i2cmcu_route[0]), .Y(n152) );
  INVX1 U696 ( .A(r_i2cslv_route[0]), .Y(n163) );
  INVX1 U697 ( .A(N262), .Y(n548) );
  OAI22AX1 U698 ( .D(n232), .C(n187), .A(n233), .B(n232), .Y(dpdm_urx) );
  OAI22X1 U699 ( .A(n146), .B(n537), .C(r_i2crout[5]), .D(n538), .Y(n232) );
  AOI22AXL U700 ( .A(n234), .B(n235), .D(n235), .C(di_gpio[0]), .Y(n233) );
  NAND3X1 U701 ( .A(N269), .B(N267), .C(N268), .Y(n235) );
  ENOX1 U702 ( .A(n236), .B(n237), .C(di_gpio[1]), .D(n236), .Y(n234) );
  NOR32XL U703 ( .B(N266), .C(N264), .A(n550), .Y(n236) );
  AOI22AXL U704 ( .A(n238), .B(di_gpio[2]), .D(n238), .C(n239), .Y(n237) );
  NOR3XL U705 ( .A(n547), .B(n549), .C(n548), .Y(n238) );
  NAND4X1 U706 ( .A(N259), .B(N260), .C(N258), .D(n240), .Y(n239) );
  INVX1 U707 ( .A(r_dpdmctl[6]), .Y(n541) );
  INVX1 U708 ( .A(r_ccctl[0]), .Y(n536) );
  NOR21XL U709 ( .B(r_do_ts[2]), .A(n66), .Y(DO_TS[2]) );
  OAI21BBX1 U710 ( .A(DI_GPIO[5]), .B(n82), .C(n170), .Y(di_gpio[5]) );
  OAI21BBX1 U711 ( .A(DI_GPIO[6]), .B(n82), .C(n169), .Y(di_gpio[6]) );
  OAI21BBX1 U712 ( .A(DI_TS), .B(n82), .C(n179), .Y(di_ts) );
  OAI221X1 U713 ( .A(r_dpdo_sel[3]), .B(n363), .C(n364), .D(n164), .E(n365), 
        .Y(n313) );
  NAND4X1 U714 ( .A(n165), .B(n164), .C(n166), .D(n366), .Y(n365) );
  AOI22X1 U715 ( .A(n383), .B(n165), .C(r_dpdo_sel[2]), .D(n384), .Y(n363) );
  AOI22X1 U716 ( .A(n369), .B(n165), .C(r_dpdo_sel[2]), .D(n370), .Y(n364) );
  OAI22X1 U717 ( .A(n377), .B(n166), .C(r_dpdo_sel[1]), .D(n378), .Y(n369) );
  AOI221XL U718 ( .A(n211), .B(di_aswk[1]), .C(n512), .D(r_ocdrv_enz), .E(n382), .Y(n377) );
  AOI221XL U719 ( .A(n211), .B(pwm_o[1]), .C(n512), .D(r_osc_stop), .E(n379), 
        .Y(n378) );
  OAI22X1 U720 ( .A(n380), .B(n139), .C(n241), .D(n381), .Y(n382) );
  AOI22X1 U721 ( .A(n406), .B(n513), .C(r_dndo_sel[3]), .D(n407), .Y(n400) );
  OAI22X1 U722 ( .A(n415), .B(n514), .C(r_dndo_sel[2]), .D(n416), .Y(n406) );
  OAI22X1 U723 ( .A(n408), .B(n514), .C(r_dndo_sel[2]), .D(n409), .Y(n407) );
  AOI222XL U724 ( .A(n412), .B(TX_DAT), .C(n515), .D(n584), .E(n519), .F(n585), 
        .Y(n416) );
  OAI22X1 U725 ( .A(r_i2crout[4]), .B(n501), .C(n148), .D(n502), .Y(n279) );
  OA22X1 U726 ( .A(n501), .B(n148), .C(n502), .D(r_i2crout[4]), .Y(CC1_DOB) );
  INVX1 U727 ( .A(sfr_intr[2]), .Y(n30) );
  NOR21XL U728 ( .B(i2c_ev_3), .A(sse_adr[7]), .Y(i2c_ev_2) );
  XNOR2XL U729 ( .A(n503), .B(r_aopt[3]), .Y(o_dodat5_2_) );
  NAND2X1 U730 ( .A(r_imp_osc), .B(di_aswk[4]), .Y(n503) );
  OAI2B11X1 U731 ( .D(r_sdischg[6]), .C(sdischg_duty), .A(n540), .B(
        r_srcctl[4]), .Y(n375) );
  OAI21BBX1 U732 ( .A(DRP_OSC), .B(n84), .C(n177), .Y(di_aswk[0]) );
  OAI21BBX1 U733 ( .A(IMP_OSC), .B(n80), .C(n177), .Y(di_aswk[4]) );
  OAI21BBX1 U734 ( .A(r_xtm[7]), .B(n554), .C(r_aopt[5]), .Y(n306) );
  OAI21X1 U735 ( .B(r_pwrctl[7]), .C(n358), .A(n359), .Y(n320) );
  OAI21X1 U736 ( .B(s0_rxdoe), .C(n146), .A(r_pwrctl[7]), .Y(n359) );
  AOI222XL U737 ( .A(r_dpdmctl[3]), .B(n360), .C(n361), .D(n146), .E(
        r_i2crout[5]), .F(n362), .Y(n358) );
  OAI22X1 U738 ( .A(slvo_sda), .B(n153), .C(mcuo_sda), .D(n149), .Y(n502) );
  OAI211X1 U739 ( .C(r_pwrctl[6]), .D(n394), .A(n395), .B(n524), .Y(n305) );
  OAI21X1 U740 ( .B(r_i2crout[5]), .C(s0_rxdoe), .A(r_pwrctl[6]), .Y(n395) );
  INVX1 U741 ( .A(fcp_oe), .Y(n524) );
  AOI222XL U742 ( .A(r_dpdmctl[1]), .B(n360), .C(r_i2crout[5]), .D(n361), .E(
        n362), .F(n146), .Y(n394) );
  OAI32X1 U743 ( .A(n508), .B(r_dpdo_sel[1]), .C(n390), .D(n391), .E(n166), 
        .Y(n383) );
  AOI22X1 U744 ( .A(r_dpdmctl[2]), .B(n584), .C(n124), .D(n542), .Y(n390) );
  AOI221XL U745 ( .A(n219), .B(n534), .C(n511), .D(n585), .E(n392), .Y(n391)
         );
  OAI22X1 U746 ( .A(n393), .B(n374), .C(n321), .D(n376), .Y(n392) );
  ENOX1 U747 ( .A(fcp_oe), .B(n404), .C(fcp_do), .D(fcp_oe), .Y(n403) );
  AOI32X1 U748 ( .A(n360), .B(n538), .C(r_dpdmctl[0]), .D(r_pwrctl[6]), .E(
        n405), .Y(n404) );
  OAI22X1 U749 ( .A(r_i2crout[5]), .B(n572), .C(n146), .D(n571), .Y(n405) );
  INVX1 U750 ( .A(r_xana_18), .Y(n139) );
  OAI22X1 U751 ( .A(n371), .B(n166), .C(r_dpdo_sel[1]), .D(n372), .Y(n370) );
  AOI221XL U752 ( .A(n219), .B(n523), .C(n511), .D(o_dodat5_2_), .E(n373), .Y(
        n371) );
  AOI222XL U753 ( .A(n511), .B(di_aswk[4]), .C(n512), .D(di_aswk[0]), .E(n219), 
        .F(r_xana_19), .Y(n372) );
  OAI22X1 U754 ( .A(n374), .B(n539), .C(n375), .D(n376), .Y(n373) );
  OAI22X1 U755 ( .A(r_dpdo_sel[1]), .B(n385), .C(n386), .D(n166), .Y(n384) );
  AOI222XL U756 ( .A(n511), .B(di_aswk[3]), .C(n211), .D(di_pro[5]), .E(n219), 
        .F(n580), .Y(n386) );
  AOI221XL U757 ( .A(n219), .B(di_pro[0]), .C(n511), .D(n581), .E(n387), .Y(
        n385) );
  OAI22X1 U758 ( .A(n388), .B(n374), .C(n389), .D(n376), .Y(n387) );
  AOI22X1 U759 ( .A(n428), .B(n514), .C(r_dndo_sel[2]), .D(n429), .Y(n426) );
  OAI22X1 U760 ( .A(r_dndo_sel[1]), .B(n430), .C(n393), .D(n517), .Y(n428) );
  OAI22X1 U761 ( .A(r_dndo_sel[1]), .B(n388), .C(n517), .D(n306), .Y(n429) );
  INVX1 U762 ( .A(r_srcctl[0]), .Y(n131) );
  INVX1 U763 ( .A(r_otpi_gate), .Y(n540) );
  OAI2B11X1 U764 ( .D(r_sdischg[5]), .C(sdischg_duty), .A(n540), .B(
        r_srcctl[1]), .Y(n425) );
  AOI21X1 U765 ( .B(RD_DET), .C(n86), .A(n594), .Y(n241) );
  NOR2X1 U766 ( .A(r_dndo_sel[0]), .B(r_dndo_sel[1]), .Y(n402) );
  NOR2X1 U767 ( .A(n517), .B(r_dndo_sel[0]), .Y(n412) );
  NAND2X1 U768 ( .A(r_dndo_sel[0]), .B(n517), .Y(n414) );
  NAND2X1 U769 ( .A(r_dpdo_sel[0]), .B(n542), .Y(n374) );
  NAND2X1 U770 ( .A(r_dpdmctl[2]), .B(n508), .Y(n376) );
  INVX1 U771 ( .A(r_pwrdn), .Y(n555) );
  NAND2X1 U772 ( .A(r_dpdo_sel[0]), .B(r_dpdmctl[2]), .Y(n380) );
  NAND2X1 U773 ( .A(r_dndo_sel[0]), .B(r_dndo_sel[1]), .Y(n411) );
  NAND2X1 U774 ( .A(r_i2cmcu_route[1]), .B(n152), .Y(n397) );
  INVX1 U775 ( .A(r_dndo_sel[1]), .Y(n517) );
  INVX1 U776 ( .A(r_dpdo_sel[0]), .Y(n508) );
  INVX1 U777 ( .A(r_dpdmctl[2]), .Y(n542) );
  INVX1 U778 ( .A(r_i2crout[4]), .Y(n148) );
  INVX1 U779 ( .A(r_vpp0v_en), .Y(n521) );
  INVX1 U780 ( .A(r_sleep), .Y(n544) );
  INVX1 U781 ( .A(r_vpp_en), .Y(n520) );
  INVX1 U782 ( .A(r_xana[12]), .Y(n141) );
  INVX1 U783 ( .A(r_srcctl[5]), .Y(n539) );
  OAI21BBX1 U784 ( .A(PMEM_Q0[7]), .B(n79), .C(n176), .Y(pmem_q0[7]) );
  OAI21BBX1 U785 ( .A(PMEM_Q1[7]), .B(n76), .C(n168), .Y(pmem_q1[7]) );
  OAI21BBX1 U786 ( .A(PMEM_Q1[1]), .B(n94), .C(n174), .Y(pmem_q1[1]) );
  OAI21BBX1 U787 ( .A(PMEM_Q0[1]), .B(n92), .C(n181), .Y(pmem_q0[1]) );
  OAI21BBX1 U788 ( .A(PMEM_Q0[2]), .B(n81), .C(n180), .Y(pmem_q0[2]) );
  OAI21BBX1 U789 ( .A(PMEM_Q1[2]), .B(n75), .C(n173), .Y(pmem_q1[2]) );
  OAI21BBX1 U790 ( .A(PMEM_Q1[3]), .B(n78), .C(n172), .Y(pmem_q1[3]) );
  OAI21BBX1 U791 ( .A(PMEM_Q0[3]), .B(n94), .C(n179), .Y(pmem_q0[3]) );
  OAI21BBX1 U792 ( .A(PMEM_Q1[5]), .B(n82), .C(n170), .Y(pmem_q1[5]) );
  OAI21BBX1 U793 ( .A(PMEM_Q0[5]), .B(n83), .C(n177), .Y(pmem_q0[5]) );
  AO22X1 U794 ( .A(n72), .B(d_dodat[14]), .C(PMEM_Q0[6]), .D(n86), .Y(
        pmem_q0[6]) );
  OAI21BBX1 U795 ( .A(PMEM_Q1[6]), .B(n74), .C(n169), .Y(pmem_q1[6]) );
  OAI21BBX1 U796 ( .A(PMEM_Q0[0]), .B(n83), .C(n182), .Y(pmem_q0[0]) );
  OAI21BBX1 U797 ( .A(PMEM_Q1[0]), .B(n80), .C(n175), .Y(pmem_q1[0]) );
  OAI21BBX1 U798 ( .A(PMEM_Q0[4]), .B(n93), .C(n178), .Y(pmem_q0[4]) );
  OAI21BBX1 U799 ( .A(PMEM_Q1[4]), .B(n92), .C(n171), .Y(pmem_q1[4]) );
  OAI21BBX1 U800 ( .A(STB_OVP), .B(n83), .C(n177), .Y(di_aswk[1]) );
  NAND2X1 U801 ( .A(r_i2cslv_route[1]), .B(n163), .Y(n396) );
  INVX1 U802 ( .A(r_i2crout[5]), .Y(n146) );
  OAI22X1 U803 ( .A(slvo_sda), .B(n396), .C(mcuo_sda), .D(n397), .Y(n361) );
  INVX1 U804 ( .A(r_dndo_sel[2]), .Y(n514) );
  INVX1 U805 ( .A(sfr_intr[3]), .Y(n31) );
  NOR2X1 U806 ( .A(r_dpdo_sel[0]), .B(n367), .Y(n366) );
  AOI32X1 U807 ( .A(n360), .B(n537), .C(r_dpdmctl[2]), .D(r_pwrctl[7]), .E(
        n368), .Y(n367) );
  OAI22X1 U808 ( .A(n146), .B(n572), .C(r_i2crout[5]), .D(n571), .Y(n368) );
  INVX1 U809 ( .A(do_opt[6]), .Y(n571) );
  INVX1 U810 ( .A(do_opt[7]), .Y(n572) );
  INVX1 U811 ( .A(r_pwrctl[6]), .Y(n538) );
  INVX1 U812 ( .A(r_pwrctl[7]), .Y(n537) );
  INVX1 U813 ( .A(r_i2c_ninc), .Y(n29) );
  OAI22X1 U814 ( .A(dp_comp), .B(n146), .C(r_i2crout[5]), .D(dm_comp), .Y(n187) );
  OAI22X1 U815 ( .A(r_i2crout[5]), .B(dp_comp), .C(dm_comp), .D(n146), .Y(n198) );
  OAI22X1 U816 ( .A(r_i2crout[4]), .B(n585), .C(n586), .D(n148), .Y(n184) );
  OAI22X1 U817 ( .A(n585), .B(n148), .C(r_i2crout[4]), .D(n586), .Y(n196) );
  INVX1 U818 ( .A(r_dpdo_sel[1]), .Y(n166) );
  INVX1 U819 ( .A(r_dndo_sel[3]), .Y(n513) );
  INVX1 U820 ( .A(r_dpdo_sel[2]), .Y(n165) );
  INVX1 U821 ( .A(r_dpdo_sel[3]), .Y(n164) );
  OAI21BBX1 U822 ( .A(t_di_gpio4), .B(n82), .C(n171), .Y(di_gpio[4]) );
  OAI21BBX1 U823 ( .A(XANAV[3]), .B(n81), .C(n172), .Y(di_xanav[3]) );
  OAI21BBX1 U824 ( .A(XANAV[2]), .B(n76), .C(n173), .Y(di_xanav[2]) );
  OAI21BBX1 U825 ( .A(XANAV[4]), .B(n81), .C(n171), .Y(di_xanav[4]) );
  NOR21XL U826 ( .B(di_tst), .A(n66), .Y(n499) );
  NOR21X2 U827 ( .B(pmem_re), .A(n90), .Y(PMEM_RE) );
  NOR21XL U828 ( .B(di_tst), .A(N595), .Y(tm_atpg) );
  NOR21XL U829 ( .B(r_do_ts[1]), .A(n66), .Y(DO_TS[1]) );
  NOR21XL U830 ( .B(r_do_ts[0]), .A(n66), .Y(DO_TS[0]) );
  NOR21XL U831 ( .B(r_pu_gpio[6]), .A(atpg_en), .Y(GPIO_PU[6]) );
  NOR21XL U832 ( .B(r_pu_gpio[5]), .A(n91), .Y(GPIO_PU[5]) );
  NOR21XL U833 ( .B(r_pu_gpio[4]), .A(n61), .Y(GPIO_PU[4]) );
  NOR21XL U836 ( .B(r_pd_gpio[3]), .A(n66), .Y(GPIO_PD[3]) );
  NOR21XL U837 ( .B(r_pd_gpio[2]), .A(n67), .Y(GPIO_PD[2]) );
  NOR21XL U838 ( .B(r_pd_gpio[1]), .A(n66), .Y(GPIO_PD[1]) );
  NOR21XL U839 ( .B(r_pd_gpio[0]), .A(n67), .Y(GPIO_PD[0]) );
  NOR21XL U840 ( .B(r_pd_gpio[6]), .A(n61), .Y(GPIO_PD[6]) );
  NOR21XL U841 ( .B(r_pd_gpio[5]), .A(n61), .Y(GPIO_PD[5]) );
  NOR21XL U842 ( .B(r_pd_gpio[4]), .A(n61), .Y(GPIO_PD[4]) );
  NOR21XL U843 ( .B(r_pu_gpio[3]), .A(n61), .Y(GPIO_PU[3]) );
  NOR21XL U844 ( .B(r_pu_gpio[2]), .A(n61), .Y(GPIO_PU[2]) );
  NOR21XL U845 ( .B(r_pu_gpio[1]), .A(n61), .Y(GPIO_PU[1]) );
  NOR21XL U846 ( .B(r_pu_gpio[0]), .A(n61), .Y(GPIO_PU[0]) );
  NOR21XL U847 ( .B(r_lt_gpi[2]), .A(n54), .Y(lt_gpi[2]) );
  NOR21XL U848 ( .B(r_lt_gpi[3]), .A(n54), .Y(lt_gpi[3]) );
  NOR21XL U849 ( .B(r_lt_gpi[1]), .A(n54), .Y(lt_gpi[1]) );
  NOR21XL U850 ( .B(r_xana[15]), .A(n62), .Y(ANA_REGX[15]) );
  NOR21XL U851 ( .B(r_xana[13]), .A(n62), .Y(ANA_REGX[13]) );
  NOR21XL U852 ( .B(r_xana[14]), .A(n62), .Y(ANA_REGX[14]) );
  NOR21XL U853 ( .B(r_regtrm[0]), .A(n90), .Y(REGTRM[0]) );
  NOR21XL U854 ( .B(r_regtrm[1]), .A(n60), .Y(REGTRM[1]) );
  NOR21XL U855 ( .B(r_regtrm[2]), .A(n59), .Y(REGTRM[2]) );
  NOR21XL U856 ( .B(r_regtrm[3]), .A(n58), .Y(REGTRM[3]) );
  NOR21XL U857 ( .B(r_regtrm[4]), .A(n57), .Y(REGTRM[4]) );
  NOR21XL U858 ( .B(r_regtrm[5]), .A(n56), .Y(REGTRM[5]) );
  NOR21XL U859 ( .B(r_regtrm[6]), .A(n56), .Y(REGTRM[6]) );
  NOR21XL U860 ( .B(r_regtrm[7]), .A(n56), .Y(REGTRM[7]) );
  NOR21XL U861 ( .B(r_regtrm[8]), .A(n56), .Y(REGTRM[8]) );
  NOR21XL U862 ( .B(r_regtrm[9]), .A(n56), .Y(REGTRM[9]) );
  NOR21XL U863 ( .B(r_regtrm[10]), .A(n91), .Y(REGTRM[10]) );
  NOR21XL U864 ( .B(r_regtrm[11]), .A(n91), .Y(REGTRM[11]) );
  NOR21XL U865 ( .B(r_regtrm[12]), .A(atpg_en), .Y(REGTRM[12]) );
  NOR21XL U866 ( .B(r_regtrm[13]), .A(n89), .Y(REGTRM[13]) );
  NOR21XL U867 ( .B(r_regtrm[14]), .A(n90), .Y(REGTRM[14]) );
  NOR21XL U868 ( .B(r_regtrm[15]), .A(n91), .Y(REGTRM[15]) );
  NOR21XL U869 ( .B(r_regtrm[16]), .A(atpg_en), .Y(REGTRM[16]) );
  NOR21XL U870 ( .B(r_regtrm[17]), .A(atpg_en), .Y(REGTRM[17]) );
  NOR21XL U871 ( .B(r_regtrm[18]), .A(n60), .Y(REGTRM[18]) );
  NOR21XL U872 ( .B(r_regtrm[19]), .A(n60), .Y(REGTRM[19]) );
  NOR21XL U873 ( .B(r_regtrm[20]), .A(n60), .Y(REGTRM[20]) );
  NOR21XL U874 ( .B(r_regtrm[21]), .A(n60), .Y(REGTRM[21]) );
  NOR21XL U875 ( .B(r_regtrm[22]), .A(n60), .Y(REGTRM[22]) );
  NOR21XL U876 ( .B(r_regtrm[23]), .A(n60), .Y(REGTRM[23]) );
  NOR21XL U877 ( .B(r_regtrm[24]), .A(n60), .Y(REGTRM[24]) );
  NOR21XL U878 ( .B(r_regtrm[25]), .A(n60), .Y(REGTRM[25]) );
  NOR21XL U879 ( .B(r_regtrm[26]), .A(n60), .Y(REGTRM[26]) );
  NOR21XL U880 ( .B(r_regtrm[27]), .A(n59), .Y(REGTRM[27]) );
  NOR21XL U881 ( .B(r_regtrm[28]), .A(n59), .Y(REGTRM[28]) );
  NOR21XL U882 ( .B(r_regtrm[29]), .A(n59), .Y(REGTRM[29]) );
  NOR21XL U883 ( .B(r_regtrm[30]), .A(n59), .Y(REGTRM[30]) );
  NOR21XL U884 ( .B(r_regtrm[31]), .A(n59), .Y(REGTRM[31]) );
  NOR21XL U885 ( .B(r_regtrm[32]), .A(n59), .Y(REGTRM[32]) );
  NOR21XL U886 ( .B(r_regtrm[33]), .A(n59), .Y(REGTRM[33]) );
  NOR21XL U887 ( .B(r_regtrm[34]), .A(n59), .Y(REGTRM[34]) );
  NOR21XL U888 ( .B(r_regtrm[35]), .A(n59), .Y(REGTRM[35]) );
  NOR21XL U889 ( .B(r_regtrm[36]), .A(n58), .Y(REGTRM[36]) );
  NOR21XL U890 ( .B(r_regtrm[37]), .A(n58), .Y(REGTRM[37]) );
  NOR21XL U891 ( .B(r_regtrm[38]), .A(n58), .Y(REGTRM[38]) );
  NOR21XL U892 ( .B(r_regtrm[39]), .A(n58), .Y(REGTRM[39]) );
  NOR21XL U893 ( .B(r_regtrm[40]), .A(n58), .Y(REGTRM[40]) );
  NOR21XL U894 ( .B(r_regtrm[41]), .A(n58), .Y(REGTRM[41]) );
  NOR21XL U895 ( .B(r_regtrm[42]), .A(n61), .Y(REGTRM[42]) );
  NOR21XL U896 ( .B(r_regtrm[43]), .A(n58), .Y(REGTRM[43]) );
  NOR21XL U897 ( .B(r_regtrm[44]), .A(n58), .Y(REGTRM[44]) );
  NOR21XL U898 ( .B(r_regtrm[45]), .A(n58), .Y(REGTRM[45]) );
  NOR21XL U899 ( .B(r_regtrm[46]), .A(n57), .Y(REGTRM[46]) );
  NOR21XL U900 ( .B(r_regtrm[47]), .A(n57), .Y(REGTRM[47]) );
  NOR21XL U901 ( .B(r_regtrm[48]), .A(n57), .Y(REGTRM[48]) );
  NOR21XL U902 ( .B(r_regtrm[49]), .A(n57), .Y(REGTRM[49]) );
  NOR21XL U903 ( .B(r_regtrm[50]), .A(n57), .Y(REGTRM[50]) );
  NOR21XL U904 ( .B(r_regtrm[51]), .A(n57), .Y(REGTRM[51]) );
  NOR21XL U905 ( .B(r_regtrm[52]), .A(n57), .Y(REGTRM[52]) );
  NOR21XL U906 ( .B(r_regtrm[53]), .A(n57), .Y(REGTRM[53]) );
  NOR21XL U907 ( .B(r_regtrm[54]), .A(n57), .Y(REGTRM[54]) );
  NOR21XL U908 ( .B(r_regtrm[55]), .A(n56), .Y(REGTRM[55]) );
  NOR21XL U909 ( .B(r_aopt[0]), .A(n61), .Y(ANAOPT[0]) );
  NOR21XL U910 ( .B(r_aopt[2]), .A(n62), .Y(ANAOPT[2]) );
  NOR21XL U911 ( .B(r_aopt[6]), .A(n62), .Y(ANAOPT[6]) );
  NOR21XL U912 ( .B(r_aopt[7]), .A(n62), .Y(ANAOPT[7]) );
  NOR21XL U913 ( .B(r_accctl[3]), .A(n65), .Y(DO_DPDN[5]) );
  NOR21XL U914 ( .B(r_cvctl[6]), .A(n65), .Y(DO_CVCTL[6]) );
  NOR21XL U915 ( .B(r_cvctl[7]), .A(n65), .Y(DO_CVCTL[7]) );
  NOR21XL U916 ( .B(r_cvctl[5]), .A(n65), .Y(DO_CVCTL[5]) );
  NOR21XL U917 ( .B(r_sdischg[7]), .A(n73), .Y(LDO3P9V) );
  NOR21XL U918 ( .B(r_ana_tm[0]), .A(n63), .Y(ANA_TM[0]) );
  NOR21XL U919 ( .B(r_ana_tm[1]), .A(n63), .Y(ANA_TM[1]) );
  NOR21XL U920 ( .B(r_ana_tm[2]), .A(n63), .Y(ANA_TM[2]) );
  NOR21XL U921 ( .B(r_ana_tm[3]), .A(n63), .Y(ANA_TM[3]) );
  NOR21XL U922 ( .B(r_cctrx[3]), .A(n64), .Y(DO_CCTRX[3]) );
  NOR21XL U923 ( .B(r_cvctl[2]), .A(n64), .Y(DO_CVCTL[2]) );
  NOR21XL U924 ( .B(r_xana_23), .A(n89), .Y(LFOSC_ENB) );
  NOR21XL U925 ( .B(r_dpdmctl[4]), .A(n65), .Y(DO_DPDN[1]) );
  NOR21XL U926 ( .B(r_dpdmctl[5]), .A(n65), .Y(DO_DPDN[2]) );
  NOR21XL U927 ( .B(r_xana[10]), .A(n62), .Y(ANA_REGX[10]) );
  NOR21XL U928 ( .B(r_xana[11]), .A(n62), .Y(ANA_REGX[11]) );
  NOR21XL U929 ( .B(r_dpdmctl[7]), .A(n65), .Y(DO_DPDN[4]) );
  NOR21XL U930 ( .B(r_accctl[4]), .A(n65), .Y(DO_DPDN[0]) );
  NOR21XL U931 ( .B(x_daclsb[2]), .A(n63), .Y(DAC1_EN) );
  NOR21XL U932 ( .B(r_cctrx[7]), .A(n64), .Y(DO_CCTRX[7]) );
  NOR21XL U933 ( .B(r_cctrx[6]), .A(n64), .Y(DO_CCTRX[6]) );
  NOR21XL U934 ( .B(r_cctrx[5]), .A(n64), .Y(DO_CCTRX[5]) );
  NOR21XL U935 ( .B(r_cctrx[4]), .A(n64), .Y(DO_CCTRX[4]) );
  NOR21XL U936 ( .B(r_xtm[0]), .A(n55), .Y(XTM[0]) );
  NOR21XL U937 ( .B(r_xtm[1]), .A(n55), .Y(XTM[1]) );
  NOR21XL U938 ( .B(r_xtm[2]), .A(n54), .Y(XTM[2]) );
  NOR21XL U939 ( .B(r_xtm[3]), .A(n54), .Y(XTM[3]) );
  NOR21XL U940 ( .B(r_cctrx[0]), .A(n64), .Y(DO_CCTRX[0]) );
  NOR21XL U941 ( .B(r_srcctl[3]), .A(n67), .Y(DO_SRCCTL[3]) );
  NOR21XL U942 ( .B(r_srcctl[2]), .A(n66), .Y(DO_SRCCTL[2]) );
  NOR21XL U943 ( .B(r_ccctl[7]), .A(n64), .Y(DO_CCCTL[7]) );
  NOR21XL U944 ( .B(r_ccctl[6]), .A(n64), .Y(DO_CCCTL[6]) );
  NOR21XL U945 ( .B(r_ccctl[4]), .A(n63), .Y(DO_CCCTL[4]) );
  NOR21XL U946 ( .B(r_ccctl[5]), .A(n64), .Y(DO_CCCTL[5]) );
  OR2X1 U947 ( .A(r_gpio_ie[0]), .B(n73), .Y(GPIO_IE[0]) );
  NOR3XL U948 ( .A(r_lt_gpi[2]), .B(r_lt_gpi[3]), .C(r_lt_gpi[1]), .Y(
        sll_223_2_A_0_) );
  NAND2X1 U949 ( .A(r_lt_gpi[0]), .B(sll_223_2_A_0_), .Y(n616) );
  NAND2X1 U950 ( .A(r_lt_gpi[0]), .B(N595), .Y(n606) );
  NAND2X1 U951 ( .A(r_lt_gpi[1]), .B(sll_223_2_A_0_), .Y(n617) );
  NAND2X1 U952 ( .A(r_lt_gpi[1]), .B(N595), .Y(n607) );
  INVX1 U953 ( .A(r_lt_gpi[3]), .Y(n577) );
  INVX1 U954 ( .A(r_lt_gpi[2]), .Y(n603) );
  NAND2X1 U955 ( .A(r_lt_gpi[2]), .B(r_lt_gpi[3]), .Y(n618) );
  NAND2X1 U956 ( .A(r_lt_gpi[2]), .B(r_lt_gpi[3]), .Y(n608) );
  NAND2X1 U957 ( .A(r_lt_gpi[2]), .B(n577), .Y(n622) );
  NAND2X1 U958 ( .A(r_lt_gpi[2]), .B(n577), .Y(n612) );
  NAND2X1 U959 ( .A(r_lt_gpi[3]), .B(n603), .Y(n624) );
  NAND2X1 U960 ( .A(r_lt_gpi[3]), .B(n603), .Y(n614) );
  OR2X1 U961 ( .A(r_gpio_ie[1]), .B(n72), .Y(GPIO_IE[1]) );
  INVX1 U962 ( .A(r_lt_gpi[0]), .Y(n604) );
  NAND2X1 U963 ( .A(di_tst), .B(n605), .Y(n327) );
  INVX1 U964 ( .A(i_rstz), .Y(n605) );
  OR2X1 U965 ( .A(r_cctrx[2]), .B(n73), .Y(DO_CCTRX[2]) );
  OR2X1 U966 ( .A(r_cctrx[1]), .B(n72), .Y(DO_CCTRX[1]) );
  AO2222XL U967 ( .A(n435), .B(di_pro[5]), .C(n436), .D(n581), .E(n143), .F(
        di_aswk[3]), .G(n440), .H(pmem_clk[0]), .Y(n441) );
  INVX1 U968 ( .A(pmem_clk[0]), .Y(n575) );
  MUX2X2 U969 ( .D0(xram_d[0]), .D1(n32), .S(n105), .Y(r_dacwdat[0]) );
  BUFX6 U970 ( .A(memaddr_c[4]), .Y(n23) );
  BUFX6 U971 ( .A(memaddr_c[2]), .Y(n24) );
  AND2X2 U972 ( .A(r_vpp0v_en), .B(ps_pwrdn), .Y(pwrdn_rst) );
  MUX2XL U973 ( .D0(xram_d[1]), .D1(n35), .S(n105), .Y(r_dacwdat[1]) );
  MUX2XL U974 ( .D0(xram_d[4]), .D1(n42), .S(n105), .Y(r_dacwdat[4]) );
  MUX2XL U975 ( .D0(xram_d[7]), .D1(n49), .S(n105), .Y(r_dacwdat[7]) );
  MUX2XL U976 ( .D0(xram_d[6]), .D1(n47), .S(n105), .Y(r_dacwdat[6]) );
  MUX2XL U977 ( .D0(xram_d[5]), .D1(n45), .S(n105), .Y(r_dacwdat[5]) );
  MUX2XL U978 ( .D0(xram_d[3]), .D1(sfr_wdat[3]), .S(n105), .Y(r_dacwdat[3])
         );
  MUX2XL U979 ( .D0(xram_d[2]), .D1(n37), .S(n2), .Y(r_dacwdat[2]) );
  BUFXL U980 ( .A(memaddr_c[1]), .Y(n27) );
  NAND21X1 U981 ( .B(wr_dacv[8]), .A(n97), .Y(n101) );
  AOI22XL U982 ( .A(n1), .B(xram_ce), .C(iram_a[4]), .D(iram_ce), .Y(n247) );
  NAND21X1 U983 ( .B(wr_dacv[12]), .A(n98), .Y(n100) );
  AOI22XL U984 ( .A(xram_a[2]), .B(xram_ce), .C(iram_a[2]), .D(iram_ce), .Y(
        n248) );
  NOR8X4 U985 ( .A(n104), .B(wr_dacv[13]), .C(n103), .D(n102), .E(n100), .F(
        r_dacwr[7]), .G(n101), .H(n99), .Y(n105) );
endmodule


module SNPS_CLOCK_GATE_HIGH_core_a0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glpwm_a0_1 ( clk, rstz, clk_base, we, wdat, r_pwm, pwm_o );
  input [7:0] wdat;
  output [7:0] r_pwm;
  input clk, rstz, clk_base, we;
  output pwm_o;
  wire   N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18, N19, N20,
         net8849, n5, n1, n2, n3, n4, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  wire   [6:0] pwmcnt;

  glreg_a0_1 u0_regpwm ( .clk(clk), .arstz(n1), .we(we), .wdat(wdat), .rdat(
        r_pwm) );
  SNPS_CLOCK_GATE_HIGH_glpwm_a0_1 clk_gate_pwmcnt_reg ( .CLK(clk_base), .EN(
        N13), .ENCLK(net8849), .TE(1'b0) );
  DFFSQX1 pwmcnt_reg_6_ ( .D(N20), .C(net8849), .XS(n2), .Q(pwmcnt[6]) );
  DFFSQX1 pwmcnt_reg_0_ ( .D(N14), .C(net8849), .XS(n1), .Q(pwmcnt[0]) );
  DFFSQX1 pwmcnt_reg_4_ ( .D(N18), .C(net8849), .XS(n2), .Q(pwmcnt[4]) );
  DFFSQX1 pwmcnt_reg_1_ ( .D(N15), .C(net8849), .XS(n1), .Q(pwmcnt[1]) );
  DFFSQX1 pwmcnt_reg_2_ ( .D(N16), .C(net8849), .XS(n2), .Q(pwmcnt[2]) );
  DFFSQX1 pwmcnt_reg_3_ ( .D(N17), .C(net8849), .XS(n2), .Q(pwmcnt[3]) );
  DFFSQX1 pwmcnt_reg_5_ ( .D(N19), .C(net8849), .XS(n2), .Q(pwmcnt[5]) );
  INVX1 U3 ( .A(n3), .Y(n1) );
  INVX1 U4 ( .A(n3), .Y(n2) );
  INVX1 U5 ( .A(rstz), .Y(n3) );
  NAND21X1 U6 ( .B(wdat[7]), .A(we), .Y(n5) );
  INVX1 U7 ( .A(n12), .Y(n25) );
  INVX1 U8 ( .A(n19), .Y(n26) );
  NAND21X1 U9 ( .B(r_pwm[7]), .A(n5), .Y(N13) );
  OAI21BBX1 U10 ( .A(N12), .B(r_pwm[7]), .C(n5), .Y(N20) );
  OAI21BBX1 U11 ( .A(N11), .B(r_pwm[7]), .C(n5), .Y(N19) );
  OAI21BBX1 U12 ( .A(N6), .B(r_pwm[7]), .C(n5), .Y(N14) );
  OAI21BBX1 U13 ( .A(N10), .B(r_pwm[7]), .C(n5), .Y(N18) );
  OAI21BBX1 U14 ( .A(N9), .B(r_pwm[7]), .C(n5), .Y(N17) );
  OAI21BBX1 U15 ( .A(N8), .B(r_pwm[7]), .C(n5), .Y(N16) );
  OAI21BBX1 U16 ( .A(N7), .B(r_pwm[7]), .C(n5), .Y(N15) );
  INVX1 U17 ( .A(pwmcnt[1]), .Y(n22) );
  INVX1 U18 ( .A(r_pwm[3]), .Y(n24) );
  INVX1 U19 ( .A(pwmcnt[5]), .Y(n21) );
  INVX1 U20 ( .A(r_pwm[2]), .Y(n23) );
  INVX1 U21 ( .A(pwmcnt[6]), .Y(n20) );
  INVX1 U22 ( .A(pwmcnt[0]), .Y(N6) );
  OR2X1 U23 ( .A(pwmcnt[1]), .B(pwmcnt[0]), .Y(n4) );
  OAI21BBX1 U24 ( .A(pwmcnt[0]), .B(pwmcnt[1]), .C(n4), .Y(N7) );
  OR2X1 U25 ( .A(n4), .B(pwmcnt[2]), .Y(n6) );
  OAI21BBX1 U26 ( .A(n4), .B(pwmcnt[2]), .C(n6), .Y(N8) );
  OR2X1 U27 ( .A(n6), .B(pwmcnt[3]), .Y(n7) );
  OAI21BBX1 U28 ( .A(n6), .B(pwmcnt[3]), .C(n7), .Y(N9) );
  OR2X1 U29 ( .A(n7), .B(pwmcnt[4]), .Y(n8) );
  OAI21BBX1 U30 ( .A(n7), .B(pwmcnt[4]), .C(n8), .Y(N10) );
  XNOR2XL U31 ( .A(n8), .B(pwmcnt[5]), .Y(N11) );
  OR2X1 U32 ( .A(pwmcnt[5]), .B(n8), .Y(n9) );
  XNOR2XL U33 ( .A(pwmcnt[6]), .B(n9), .Y(N12) );
  NOR2X1 U34 ( .A(n20), .B(r_pwm[6]), .Y(n19) );
  OR2X1 U35 ( .A(r_pwm[5]), .B(n21), .Y(n11) );
  NOR32XL U36 ( .B(r_pwm[4]), .C(n11), .A(pwmcnt[4]), .Y(n10) );
  AOI221XL U37 ( .A(r_pwm[6]), .B(n20), .C(r_pwm[5]), .D(n21), .E(n10), .Y(n18) );
  OAI2B11X1 U38 ( .D(pwmcnt[4]), .C(r_pwm[4]), .A(n11), .B(n26), .Y(n17) );
  AND2X1 U39 ( .A(pwmcnt[3]), .B(n24), .Y(n15) );
  OAI32X1 U40 ( .A(n23), .B(pwmcnt[2]), .C(n15), .D(pwmcnt[3]), .E(n24), .Y(
        n12) );
  AOI21BBXL U41 ( .B(n22), .C(r_pwm[1]), .A(pwmcnt[0]), .Y(n13) );
  AOI221XL U42 ( .A(r_pwm[1]), .B(n22), .C(n13), .D(r_pwm[0]), .E(n12), .Y(n14) );
  GEN2XL U43 ( .D(pwmcnt[2]), .E(n23), .C(n15), .B(n25), .A(n14), .Y(n16) );
  OAI22X1 U44 ( .A(n19), .B(n18), .C(n17), .D(n16), .Y(pwm_o) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glpwm_a0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_1 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net8867;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_1 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net8867), .TE(1'b0) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net8867), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net8867), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net8867), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net8867), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net8867), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net8867), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net8867), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net8867), .XR(arstz), .Q(rdat[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glpwm_a0_0 ( clk, rstz, clk_base, we, wdat, r_pwm, pwm_o );
  input [7:0] wdat;
  output [7:0] r_pwm;
  input clk, rstz, clk_base, we;
  output pwm_o;
  wire   N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18, N19, N20,
         net8885, n5, n1, n2, n3, n4, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  wire   [6:0] pwmcnt;

  glreg_a0_0 u0_regpwm ( .clk(clk), .arstz(n1), .we(we), .wdat(wdat), .rdat(
        r_pwm) );
  SNPS_CLOCK_GATE_HIGH_glpwm_a0_0 clk_gate_pwmcnt_reg ( .CLK(clk_base), .EN(
        N13), .ENCLK(net8885), .TE(1'b0) );
  DFFSQX1 pwmcnt_reg_6_ ( .D(N20), .C(net8885), .XS(n2), .Q(pwmcnt[6]) );
  DFFSQX1 pwmcnt_reg_0_ ( .D(N14), .C(net8885), .XS(n1), .Q(pwmcnt[0]) );
  DFFSQX1 pwmcnt_reg_4_ ( .D(N18), .C(net8885), .XS(n2), .Q(pwmcnt[4]) );
  DFFSQX1 pwmcnt_reg_1_ ( .D(N15), .C(net8885), .XS(n1), .Q(pwmcnt[1]) );
  DFFSQX1 pwmcnt_reg_2_ ( .D(N16), .C(net8885), .XS(n2), .Q(pwmcnt[2]) );
  DFFSQX1 pwmcnt_reg_3_ ( .D(N17), .C(net8885), .XS(n2), .Q(pwmcnt[3]) );
  DFFSQX1 pwmcnt_reg_5_ ( .D(N19), .C(net8885), .XS(n2), .Q(pwmcnt[5]) );
  INVX1 U3 ( .A(n3), .Y(n1) );
  INVX1 U4 ( .A(n3), .Y(n2) );
  INVX1 U5 ( .A(rstz), .Y(n3) );
  NAND21X1 U6 ( .B(wdat[7]), .A(we), .Y(n5) );
  INVX1 U7 ( .A(n12), .Y(n25) );
  INVX1 U8 ( .A(n19), .Y(n26) );
  NAND21X1 U9 ( .B(r_pwm[7]), .A(n5), .Y(N13) );
  OAI21BBX1 U10 ( .A(N12), .B(r_pwm[7]), .C(n5), .Y(N20) );
  OAI21BBX1 U11 ( .A(N11), .B(r_pwm[7]), .C(n5), .Y(N19) );
  OAI21BBX1 U12 ( .A(N6), .B(r_pwm[7]), .C(n5), .Y(N14) );
  OAI21BBX1 U13 ( .A(N10), .B(r_pwm[7]), .C(n5), .Y(N18) );
  OAI21BBX1 U14 ( .A(N9), .B(r_pwm[7]), .C(n5), .Y(N17) );
  OAI21BBX1 U15 ( .A(N8), .B(r_pwm[7]), .C(n5), .Y(N16) );
  OAI21BBX1 U16 ( .A(N7), .B(r_pwm[7]), .C(n5), .Y(N15) );
  INVX1 U17 ( .A(pwmcnt[1]), .Y(n22) );
  INVX1 U18 ( .A(r_pwm[3]), .Y(n24) );
  INVX1 U19 ( .A(pwmcnt[5]), .Y(n21) );
  INVX1 U20 ( .A(r_pwm[2]), .Y(n23) );
  INVX1 U21 ( .A(pwmcnt[6]), .Y(n20) );
  INVX1 U22 ( .A(pwmcnt[0]), .Y(N6) );
  OR2X1 U23 ( .A(pwmcnt[1]), .B(pwmcnt[0]), .Y(n4) );
  OAI21BBX1 U24 ( .A(pwmcnt[0]), .B(pwmcnt[1]), .C(n4), .Y(N7) );
  OR2X1 U25 ( .A(n4), .B(pwmcnt[2]), .Y(n6) );
  OAI21BBX1 U26 ( .A(n4), .B(pwmcnt[2]), .C(n6), .Y(N8) );
  OR2X1 U27 ( .A(n6), .B(pwmcnt[3]), .Y(n7) );
  OAI21BBX1 U28 ( .A(n6), .B(pwmcnt[3]), .C(n7), .Y(N9) );
  OR2X1 U29 ( .A(n7), .B(pwmcnt[4]), .Y(n8) );
  OAI21BBX1 U30 ( .A(n7), .B(pwmcnt[4]), .C(n8), .Y(N10) );
  XNOR2XL U31 ( .A(n8), .B(pwmcnt[5]), .Y(N11) );
  OR2X1 U32 ( .A(pwmcnt[5]), .B(n8), .Y(n9) );
  XNOR2XL U33 ( .A(pwmcnt[6]), .B(n9), .Y(N12) );
  NOR2X1 U34 ( .A(n20), .B(r_pwm[6]), .Y(n19) );
  OR2X1 U35 ( .A(r_pwm[5]), .B(n21), .Y(n11) );
  NOR32XL U36 ( .B(r_pwm[4]), .C(n11), .A(pwmcnt[4]), .Y(n10) );
  AOI221XL U37 ( .A(r_pwm[6]), .B(n20), .C(r_pwm[5]), .D(n21), .E(n10), .Y(n18) );
  OAI2B11X1 U38 ( .D(pwmcnt[4]), .C(r_pwm[4]), .A(n11), .B(n26), .Y(n17) );
  AND2X1 U39 ( .A(pwmcnt[3]), .B(n24), .Y(n15) );
  OAI32X1 U40 ( .A(n23), .B(pwmcnt[2]), .C(n15), .D(pwmcnt[3]), .E(n24), .Y(
        n12) );
  AOI21BBXL U41 ( .B(n22), .C(r_pwm[1]), .A(pwmcnt[0]), .Y(n13) );
  AOI221XL U42 ( .A(r_pwm[1]), .B(n22), .C(n13), .D(r_pwm[0]), .E(n12), .Y(n14) );
  GEN2XL U43 ( .D(pwmcnt[2]), .E(n23), .C(n15), .B(n25), .A(n14), .Y(n16) );
  OAI22X1 U44 ( .A(n19), .B(n18), .C(n17), .D(n16), .Y(pwm_o) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glpwm_a0_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_0 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net8903;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_0 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net8903), .TE(1'b0) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net8903), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net8903), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net8903), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net8903), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net8903), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net8903), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net8903), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net8903), .XR(arstz), .Q(rdat[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module divclk_a0 ( mclk, srstz, atpg_en, clk_1500k, clk_500k, clk_100k, 
        clk_50k, clk_500, divff_8, divff_5 );
  input mclk, srstz, atpg_en;
  output clk_1500k, clk_500k, clk_100k, clk_50k, clk_500, divff_8, divff_5;
  wire   div100k_2, N11, N12, N17, N18, N24, N25, N26, N33, N34, N35, N36, N37,
         N38, N39, N40, N41, N42, N43, N44, N45, N46, n4, n5, n6, n7, n8, n9,
         n10, n1, n2, n3, n11, n12, n13;
  wire   [1:0] div8;
  wire   [1:0] div500k_5;
  wire   [1:0] div1p5m_3;
  wire   [6:0] div50k_100;

  CLKDLX1 U0_D1P5M_ICG ( .CK(mclk), .E(n7), .SE(atpg_en), .ECK(clk_1500k) );
  CLKDLX1 U0_D500K_ICG ( .CK(clk_1500k), .E(n8), .SE(atpg_en), .ECK(clk_500k)
         );
  CLKDLX1 U0_D100K_ICG ( .CK(clk_500k), .E(n9), .SE(atpg_en), .ECK(clk_100k)
         );
  CLKDLX1 U0_D50K_ICG ( .CK(clk_100k), .E(div100k_2), .SE(atpg_en), .ECK(
        clk_50k) );
  CLKDLX1 U0_D0P5K_ICG ( .CK(clk_50k), .E(n10), .SE(atpg_en), .ECK(clk_500) );
  divclk_a0_DW01_inc_0 add_48 ( .A(div50k_100), .SUM({N39, N38, N37, N36, N35, 
        N34, N33}) );
  DFFRQX1 div100k_2_reg ( .D(n13), .C(clk_100k), .XR(n1), .Q(div100k_2) );
  DFFRQX1 div50k_100_reg_6_ ( .D(N46), .C(clk_50k), .XR(n2), .Q(div50k_100[6])
         );
  DFFRQX1 div50k_100_reg_5_ ( .D(N45), .C(clk_50k), .XR(n2), .Q(div50k_100[5])
         );
  DFFRQX1 div50k_100_reg_4_ ( .D(N44), .C(clk_50k), .XR(n2), .Q(div50k_100[4])
         );
  DFFRQX1 div1p5m_3_reg_1_ ( .D(N18), .C(clk_1500k), .XR(n1), .Q(div1p5m_3[1])
         );
  DFFRQX1 div1p5m_3_reg_0_ ( .D(N17), .C(clk_1500k), .XR(n1), .Q(div1p5m_3[0])
         );
  DFFRQX1 div8_reg_1_ ( .D(N11), .C(mclk), .XR(n1), .Q(div8[1]) );
  DFFRQX1 div8_reg_0_ ( .D(n11), .C(mclk), .XR(n1), .Q(div8[0]) );
  DFFRQX1 div50k_100_reg_1_ ( .D(N41), .C(clk_50k), .XR(n2), .Q(div50k_100[1])
         );
  DFFRQX1 div50k_100_reg_0_ ( .D(N40), .C(clk_50k), .XR(n1), .Q(div50k_100[0])
         );
  DFFRQX1 div50k_100_reg_3_ ( .D(N43), .C(clk_50k), .XR(n2), .Q(div50k_100[3])
         );
  DFFRQX1 div50k_100_reg_2_ ( .D(N42), .C(clk_50k), .XR(n2), .Q(div50k_100[2])
         );
  DFFRQX1 div500k_5_reg_0_ ( .D(N24), .C(clk_500k), .XR(n1), .Q(div500k_5[0])
         );
  DFFRQX1 div500k_5_reg_1_ ( .D(N25), .C(clk_500k), .XR(n1), .Q(div500k_5[1])
         );
  DFFRQX1 div8_reg_2_ ( .D(N12), .C(mclk), .XR(n1), .Q(divff_8) );
  DFFRQX1 div500k_5_reg_2_ ( .D(N26), .C(clk_500k), .XR(n1), .Q(divff_5) );
  INVX1 U3 ( .A(n3), .Y(n1) );
  INVX1 U4 ( .A(n3), .Y(n2) );
  INVX1 U5 ( .A(srstz), .Y(n3) );
  NOR21XL U6 ( .B(N38), .A(n10), .Y(N45) );
  NOR21XL U7 ( .B(N37), .A(n10), .Y(N44) );
  NOR21XL U8 ( .B(N36), .A(n10), .Y(N43) );
  NOR21XL U9 ( .B(N35), .A(n10), .Y(N42) );
  NOR21XL U10 ( .B(N34), .A(n10), .Y(N41) );
  NOR21XL U11 ( .B(N39), .A(n10), .Y(N46) );
  NOR21XL U12 ( .B(N33), .A(n10), .Y(N40) );
  XNOR2XL U13 ( .A(n12), .B(div500k_5[0]), .Y(N25) );
  AND4X1 U14 ( .A(div50k_100[5]), .B(div50k_100[1]), .C(div50k_100[6]), .D(n5), 
        .Y(n10) );
  NOR41XL U15 ( .D(div50k_100[0]), .A(div50k_100[4]), .B(div50k_100[3]), .C(
        div50k_100[2]), .Y(n5) );
  ENOX1 U16 ( .A(divff_5), .B(n4), .C(N25), .D(divff_5), .Y(N26) );
  INVX1 U17 ( .A(div500k_5[1]), .Y(n12) );
  NOR32XL U18 ( .B(divff_5), .C(n4), .A(N25), .Y(n9) );
  NOR32XL U19 ( .B(divff_8), .C(n11), .A(div8[1]), .Y(n7) );
  NOR21XL U20 ( .B(div1p5m_3[0]), .A(div1p5m_3[1]), .Y(N18) );
  NOR21XL U21 ( .B(div1p5m_3[1]), .A(div1p5m_3[0]), .Y(n8) );
  XNOR2XL U22 ( .A(divff_8), .B(n6), .Y(N12) );
  NAND2X1 U23 ( .A(div8[1]), .B(div8[0]), .Y(n6) );
  XNOR2XL U24 ( .A(n11), .B(div8[1]), .Y(N11) );
  AOI21X1 U25 ( .B(divff_5), .C(n12), .A(div500k_5[0]), .Y(N24) );
  INVX1 U26 ( .A(div8[0]), .Y(n11) );
  NOR2X1 U27 ( .A(div1p5m_3[1]), .B(div1p5m_3[0]), .Y(N17) );
  NAND2X1 U28 ( .A(div500k_5[1]), .B(div500k_5[0]), .Y(n4) );
  INVX1 U29 ( .A(div100k_2), .Y(n13) );
endmodule


module divclk_a0_DW01_inc_0 ( A, SUM );
  input [6:0] A;
  output [6:0] SUM;

  wire   [6:2] carry;

  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  XOR2X1 U1 ( .A(carry[6]), .B(A[6]), .Y(SUM[6]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module srambist_a0 ( clk, srstz, reg_hit, reg_w, reg_r, reg_wdat, iram_rdat, 
        xram_rdat, bist_en, bist_xram, bist_wr, bist_adr, bist_wdat, o_bistctl, 
        o_bistdat );
  input [1:0] reg_hit;
  input [7:0] reg_wdat;
  input [7:0] iram_rdat;
  input [7:0] xram_rdat;
  output [10:0] bist_adr;
  output [7:0] bist_wdat;
  output [6:0] o_bistctl;
  output [7:0] o_bistdat;
  input clk, srstz, reg_w, reg_r;
  output bist_en, bist_xram, bist_wr;
  wire   we_1_, bistctl_re, N21, busy_dly, N53, N54, N55, N56, N57, N58, N59,
         N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N73,
         N74, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97,
         r_bistfault, upd_fault, wd_fault, net8921, n30, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n3, n4, n5, n6, n7, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n31, n32, n33, n34, n93, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123;
  wire   [1:0] rw_sta;

  glreg_WIDTH1_0 u0_bistfault ( .clk(clk), .arstz(n11), .we(upd_fault), .wdat(
        wd_fault), .rdat(o_bistctl[3]) );
  glreg_WIDTH5_1 u0_bistctl ( .clk(clk), .arstz(n11), .we(n30), .wdat({
        reg_wdat[6:4], reg_wdat[2:1]}), .rdat({o_bistctl[6:4], o_bistctl[2:1]}) );
  glreg_a0_6 u0_bistdat ( .clk(clk), .arstz(n10), .we(we_1_), .wdat(reg_wdat), 
        .rdat(o_bistdat) );
  SNPS_CLOCK_GATE_HIGH_srambist_a0 clk_gate_adr_reg ( .CLK(clk), .EN(N86), 
        .ENCLK(net8921), .TE(1'b0) );
  srambist_a0_DW01_inc_0 add_65 ( .A(bist_adr), .SUM({N74, N73, N72, N71, N70, 
        N69, N68, N67, N66, N65, N64}) );
  DFFQX1 busy_dly_reg ( .D(o_bistctl[0]), .C(clk), .Q(busy_dly) );
  DFFQX1 r_bistfault_reg ( .D(n110), .C(clk), .Q(r_bistfault) );
  DFFRQX1 bistctl_re_reg ( .D(N21), .C(clk), .XR(n11), .Q(bistctl_re) );
  DFFQX1 rw_sta_reg_0_ ( .D(n111), .C(clk), .Q(rw_sta[0]) );
  DFFQX1 rw_sta_reg_1_ ( .D(n93), .C(clk), .Q(rw_sta[1]) );
  DFFQX1 adr_reg_9_ ( .D(N96), .C(net8921), .Q(bist_adr[9]) );
  DFFQX1 adr_reg_10_ ( .D(N97), .C(net8921), .Q(bist_adr[10]) );
  DFFQX1 adr_reg_8_ ( .D(N95), .C(net8921), .Q(bist_adr[8]) );
  DFFQX1 adr_reg_6_ ( .D(N93), .C(net8921), .Q(bist_adr[6]) );
  DFFQX1 adr_reg_7_ ( .D(N94), .C(net8921), .Q(bist_adr[7]) );
  DFFQX1 adr_reg_3_ ( .D(N90), .C(net8921), .Q(bist_adr[3]) );
  DFFQX1 adr_reg_2_ ( .D(N89), .C(net8921), .Q(bist_adr[2]) );
  DFFQX1 adr_reg_1_ ( .D(N88), .C(net8921), .Q(bist_adr[1]) );
  DFFQX1 adr_reg_0_ ( .D(N87), .C(net8921), .Q(bist_adr[0]) );
  DFFQX1 adr_reg_4_ ( .D(N91), .C(net8921), .Q(bist_adr[4]) );
  DFFQX1 adr_reg_5_ ( .D(N92), .C(net8921), .Q(bist_adr[5]) );
  INVX1 U3 ( .A(1'b1), .Y(bist_xram) );
  OR2X1 U5 ( .A(n107), .B(n106), .Y(n3) );
  INVXL U6 ( .A(n3), .Y(n4) );
  INVXL U7 ( .A(n3), .Y(n5) );
  INVXL U8 ( .A(n91), .Y(n6) );
  INVXL U9 ( .A(n6), .Y(n7) );
  INVX1 U10 ( .A(n115), .Y(bist_en) );
  INVX1 U11 ( .A(n13), .Y(n11) );
  INVX1 U12 ( .A(n13), .Y(n12) );
  INVX1 U13 ( .A(n13), .Y(n10) );
  INVX1 U14 ( .A(srstz), .Y(n13) );
  INVX1 U15 ( .A(n108), .Y(n30) );
  NAND2X1 U16 ( .A(reg_hit[0]), .B(reg_w), .Y(n108) );
  AND2X1 U17 ( .A(reg_w), .B(reg_hit[1]), .Y(we_1_) );
  XOR2X1 U18 ( .A(bist_wdat[2]), .B(iram_rdat[2]), .Y(n48) );
  XNOR2XL U19 ( .A(bist_wdat[4]), .B(n122), .Y(n44) );
  INVX1 U20 ( .A(iram_rdat[4]), .Y(n122) );
  INVX1 U21 ( .A(iram_rdat[6]), .Y(n120) );
  INVX1 U22 ( .A(iram_rdat[5]), .Y(n121) );
  INVX1 U23 ( .A(n86), .Y(n27) );
  INVX1 U24 ( .A(n76), .Y(n113) );
  INVX1 U25 ( .A(n57), .Y(n31) );
  NAND21X1 U26 ( .B(n107), .A(n106), .Y(n91) );
  NOR2X1 U27 ( .A(n105), .B(n106), .Y(n94) );
  NAND3X1 U28 ( .A(n105), .B(n11), .C(n107), .Y(N86) );
  AND2X1 U29 ( .A(reg_r), .B(reg_hit[0]), .Y(N21) );
  NAND21X1 U30 ( .B(n89), .A(n23), .Y(n84) );
  NAND2X1 U31 ( .A(n87), .B(n84), .Y(bist_wdat[0]) );
  OAI22X1 U32 ( .A(n23), .B(n86), .C(n27), .D(n84), .Y(bist_wdat[4]) );
  NAND2X1 U33 ( .A(n28), .B(n83), .Y(n86) );
  XNOR2XL U34 ( .A(n23), .B(n90), .Y(bist_wdat[1]) );
  AOI21X1 U35 ( .B(n86), .C(n28), .A(n89), .Y(n90) );
  NOR4XL U36 ( .A(n65), .B(n66), .C(n67), .D(n68), .Y(n49) );
  XNOR2XL U37 ( .A(n73), .B(n121), .Y(n65) );
  XNOR2XL U38 ( .A(n24), .B(iram_rdat[7]), .Y(n66) );
  XNOR2XL U39 ( .A(n71), .B(n72), .Y(n67) );
  INVX1 U40 ( .A(n85), .Y(n28) );
  XNOR2XL U41 ( .A(n23), .B(n88), .Y(bist_wdat[2]) );
  AOI21X1 U42 ( .B(n86), .C(n83), .A(n89), .Y(n88) );
  XNOR2XL U43 ( .A(n56), .B(n122), .Y(n55) );
  OAI22X1 U44 ( .A(n24), .B(n57), .C(n31), .D(n25), .Y(n56) );
  OAI22X1 U45 ( .A(n84), .B(n28), .C(n85), .D(n23), .Y(bist_wdat[5]) );
  OAI221X1 U46 ( .A(n84), .B(n86), .C(n27), .D(n23), .E(n87), .Y(bist_wdat[3])
         );
  INVX1 U47 ( .A(iram_rdat[0]), .Y(n123) );
  NOR4XL U48 ( .A(n41), .B(n42), .C(n43), .D(n44), .Y(n39) );
  XNOR2XL U49 ( .A(bist_wdat[0]), .B(n123), .Y(n41) );
  XOR2X1 U50 ( .A(bist_wdat[3]), .B(iram_rdat[3]), .Y(n43) );
  XNOR2XL U51 ( .A(bist_wdat[6]), .B(n120), .Y(n42) );
  NOR4XL U52 ( .A(n45), .B(n46), .C(n47), .D(n48), .Y(n38) );
  XNOR2XL U53 ( .A(bist_wdat[5]), .B(n121), .Y(n45) );
  XOR2X1 U54 ( .A(bist_wdat[1]), .B(iram_rdat[1]), .Y(n47) );
  XNOR2XL U55 ( .A(n23), .B(iram_rdat[7]), .Y(n46) );
  NOR4XL U56 ( .A(n52), .B(n53), .C(n54), .D(n55), .Y(n50) );
  XNOR2XL U57 ( .A(n63), .B(n123), .Y(n52) );
  XNOR2XL U58 ( .A(n61), .B(n120), .Y(n53) );
  XNOR2XL U59 ( .A(iram_rdat[3]), .B(n58), .Y(n54) );
  NOR2X1 U60 ( .A(n51), .B(n115), .Y(bist_wr) );
  INVX1 U61 ( .A(o_bistctl[0]), .Y(n115) );
  OAI21X1 U62 ( .B(n115), .C(n77), .A(n12), .Y(n76) );
  NOR2X1 U63 ( .A(n114), .B(n118), .Y(n77) );
  NAND2X1 U64 ( .A(n32), .B(n62), .Y(n57) );
  OAI22X1 U65 ( .A(n25), .B(n32), .C(n74), .D(n24), .Y(n73) );
  AOI21X1 U66 ( .B(n57), .C(n32), .A(n64), .Y(n71) );
  NAND3X1 U67 ( .A(n114), .B(n118), .C(n11), .Y(n40) );
  INVX1 U68 ( .A(n59), .Y(n25) );
  INVX1 U69 ( .A(n74), .Y(n32) );
  OAI22X1 U70 ( .A(n114), .B(n76), .C(n113), .D(n40), .Y(n111) );
  NAND2X1 U71 ( .A(n60), .B(n25), .Y(n63) );
  NAND42X1 U72 ( .C(o_bistdat[6]), .D(n108), .A(reg_wdat[0]), .B(o_bistdat[7]), 
        .Y(n105) );
  AOI22AXL U73 ( .A(o_bistctl[1]), .B(n108), .D(n108), .C(reg_wdat[1]), .Y(
        n106) );
  OAI2B11X1 U74 ( .D(N74), .C(n7), .A(n10), .B(n92), .Y(N97) );
  AOI21X1 U75 ( .B(N63), .C(n4), .A(n94), .Y(n92) );
  OAI2B11X1 U76 ( .D(N64), .C(n91), .A(n12), .B(n104), .Y(N87) );
  AOI21X1 U77 ( .B(N53), .C(n4), .A(n94), .Y(n104) );
  OAI2B11X1 U78 ( .D(N72), .C(n91), .A(n10), .B(n96), .Y(N95) );
  AOI21X1 U79 ( .B(N61), .C(n5), .A(n94), .Y(n96) );
  OAI2B11X1 U80 ( .D(N71), .C(n7), .A(n12), .B(n97), .Y(N94) );
  AOI21X1 U81 ( .B(N60), .C(n4), .A(n94), .Y(n97) );
  OAI2B11X1 U82 ( .D(N70), .C(n91), .A(n12), .B(n98), .Y(N93) );
  AOI21X1 U83 ( .B(N59), .C(n5), .A(n94), .Y(n98) );
  OAI2B11X1 U84 ( .D(N69), .C(n7), .A(n12), .B(n99), .Y(N92) );
  AOI21X1 U85 ( .B(N58), .C(n4), .A(n94), .Y(n99) );
  OAI2B11X1 U86 ( .D(N68), .C(n91), .A(n12), .B(n100), .Y(N91) );
  AOI21X1 U87 ( .B(N57), .C(n5), .A(n94), .Y(n100) );
  OAI2B11X1 U88 ( .D(N67), .C(n7), .A(n12), .B(n101), .Y(N90) );
  AOI21X1 U89 ( .B(N56), .C(n4), .A(n94), .Y(n101) );
  OAI2B11X1 U90 ( .D(N66), .C(n91), .A(n12), .B(n102), .Y(N89) );
  AOI21X1 U91 ( .B(N55), .C(n5), .A(n94), .Y(n102) );
  OAI2B11X1 U92 ( .D(N65), .C(n7), .A(n12), .B(n103), .Y(N88) );
  AOI21X1 U93 ( .B(N54), .C(n5), .A(n94), .Y(n103) );
  NAND2X1 U94 ( .A(n109), .B(n105), .Y(n107) );
  OAI32X1 U95 ( .A(n118), .B(rw_sta[0]), .C(n34), .D(o_bistctl[2]), .E(n51), 
        .Y(n109) );
  INVX1 U96 ( .A(o_bistctl[2]), .Y(n34) );
  OAI2B11X1 U97 ( .D(N73), .C(n7), .A(srstz), .B(n95), .Y(N96) );
  NAND2X1 U98 ( .A(N62), .B(n4), .Y(n95) );
  AND4X1 U99 ( .A(bist_adr[8]), .B(bist_adr[6]), .C(bist_adr[7]), .D(
        bist_adr[5]), .Y(n80) );
  NAND3X1 U100 ( .A(bist_adr[10]), .B(n78), .C(bist_adr[9]), .Y(o_bistctl[0])
         );
  AO44X1 U101 ( .A(bist_adr[4]), .B(bist_adr[3]), .C(n79), .D(n80), .E(n116), 
        .F(n117), .G(n81), .H(n82), .Y(n78) );
  INVX1 U102 ( .A(bist_adr[4]), .Y(n116) );
  INVX1 U103 ( .A(bist_adr[5]), .Y(n117) );
  AND3X1 U104 ( .A(bist_adr[2]), .B(bist_adr[0]), .C(bist_adr[1]), .Y(n79) );
  NOR4XL U105 ( .A(bist_adr[3]), .B(bist_adr[2]), .C(bist_adr[1]), .D(
        bist_adr[0]), .Y(n82) );
  NOR3XL U106 ( .A(bist_adr[6]), .B(bist_adr[8]), .C(bist_adr[7]), .Y(n81) );
  INVX1 U107 ( .A(o_bistdat[5]), .Y(n23) );
  NOR2X1 U108 ( .A(o_bistdat[3]), .B(o_bistdat[2]), .Y(n89) );
  NAND2X1 U109 ( .A(o_bistdat[5]), .B(n89), .Y(n87) );
  BUFX3 U110 ( .A(o_bistdat[5]), .Y(bist_wdat[7]) );
  XNOR2XL U111 ( .A(n69), .B(n70), .Y(n68) );
  AOI21X1 U112 ( .B(n57), .C(n62), .A(n64), .Y(n69) );
  XNOR2XL U113 ( .A(o_bistdat[4]), .B(iram_rdat[2]), .Y(n70) );
  NOR2X1 U114 ( .A(n29), .B(o_bistdat[2]), .Y(n85) );
  OAI31XL U115 ( .A(n119), .B(bistctl_re), .C(n13), .D(n35), .Y(n110) );
  AOI33X1 U116 ( .A(n12), .B(n112), .C(n36), .D(o_bistctl[2]), .E(busy_dly), 
        .F(n37), .Y(n35) );
  AOI211X1 U117 ( .C(n38), .D(n39), .A(n40), .B(bistctl_re), .Y(n37) );
  AOI21X1 U118 ( .B(n49), .C(n50), .A(n51), .Y(n36) );
  NAND2X1 U119 ( .A(o_bistdat[2]), .B(n29), .Y(n83) );
  INVX1 U120 ( .A(o_bistdat[3]), .Y(n29) );
  XNOR2XL U121 ( .A(o_bistdat[4]), .B(iram_rdat[1]), .Y(n72) );
  ENOX1 U122 ( .A(n83), .B(n84), .C(n83), .D(o_bistdat[5]), .Y(bist_wdat[6])
         );
  NOR2X1 U123 ( .A(n33), .B(o_bistdat[0]), .Y(n74) );
  NOR2X1 U124 ( .A(n64), .B(o_bistdat[4]), .Y(n59) );
  NAND2X1 U125 ( .A(o_bistdat[4]), .B(n64), .Y(n60) );
  NOR2X1 U126 ( .A(o_bistdat[1]), .B(o_bistdat[0]), .Y(n64) );
  AOI221XL U127 ( .A(o_bistdat[4]), .B(n57), .C(n31), .D(n59), .E(n26), .Y(n58) );
  INVX1 U128 ( .A(n60), .Y(n26) );
  ENOX1 U129 ( .A(n62), .B(n25), .C(n62), .D(o_bistdat[4]), .Y(n61) );
  INVX1 U130 ( .A(rw_sta[1]), .Y(n118) );
  NAND2X1 U131 ( .A(o_bistdat[0]), .B(n33), .Y(n62) );
  NAND2X1 U132 ( .A(rw_sta[0]), .B(n118), .Y(n51) );
  INVX1 U133 ( .A(o_bistdat[1]), .Y(n33) );
  INVX1 U134 ( .A(n75), .Y(n93) );
  AOI32X1 U135 ( .A(bist_wr), .B(n11), .C(o_bistctl[2]), .D(rw_sta[1]), .E(
        n113), .Y(n75) );
  INVX1 U136 ( .A(o_bistdat[4]), .Y(n24) );
  INVX1 U137 ( .A(rw_sta[0]), .Y(n114) );
  INVX1 U138 ( .A(bistctl_re), .Y(n112) );
  NOR2X1 U139 ( .A(bistctl_re), .B(n119), .Y(wd_fault) );
  NAND2X1 U140 ( .A(n119), .B(n112), .Y(upd_fault) );
  INVX1 U141 ( .A(r_bistfault), .Y(n119) );
  INVX1 U142 ( .A(bist_adr[0]), .Y(N53) );
  OR2X1 U143 ( .A(bist_adr[1]), .B(bist_adr[0]), .Y(n15) );
  OR2X1 U144 ( .A(n15), .B(bist_adr[2]), .Y(n16) );
  OR2X1 U145 ( .A(n16), .B(bist_adr[3]), .Y(n17) );
  OR2X1 U146 ( .A(n17), .B(bist_adr[4]), .Y(n18) );
  OR2X1 U147 ( .A(n18), .B(bist_adr[5]), .Y(n19) );
  OR2X1 U148 ( .A(n19), .B(bist_adr[6]), .Y(n20) );
  OR2X1 U149 ( .A(n20), .B(bist_adr[7]), .Y(n21) );
  OR2X1 U150 ( .A(n21), .B(bist_adr[8]), .Y(n22) );
  OR2X1 U151 ( .A(bist_adr[9]), .B(n22), .Y(n14) );
  XNOR2XL U152 ( .A(bist_adr[10]), .B(n14), .Y(N63) );
  OAI21BBX1 U153 ( .A(bist_adr[0]), .B(bist_adr[1]), .C(n15), .Y(N54) );
  OAI21BBX1 U154 ( .A(n15), .B(bist_adr[2]), .C(n16), .Y(N55) );
  OAI21BBX1 U155 ( .A(n16), .B(bist_adr[3]), .C(n17), .Y(N56) );
  OAI21BBX1 U156 ( .A(n17), .B(bist_adr[4]), .C(n18), .Y(N57) );
  OAI21BBX1 U157 ( .A(n18), .B(bist_adr[5]), .C(n19), .Y(N58) );
  OAI21BBX1 U158 ( .A(n19), .B(bist_adr[6]), .C(n20), .Y(N59) );
  OAI21BBX1 U159 ( .A(n20), .B(bist_adr[7]), .C(n21), .Y(N60) );
  OAI21BBX1 U160 ( .A(n21), .B(bist_adr[8]), .C(n22), .Y(N61) );
  XNOR2XL U161 ( .A(n22), .B(bist_adr[9]), .Y(N62) );
endmodule


module srambist_a0_DW01_inc_0 ( A, SUM );
  input [10:0] A;
  output [10:0] SUM;

  wire   [10:2] carry;

  HAD1X1 U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .SO(SUM[9]) );
  HAD1X1 U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .SO(SUM[8]) );
  HAD1X1 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .SO(SUM[7]) );
  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  XOR2X1 U1 ( .A(carry[10]), .B(A[10]), .Y(SUM[10]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_srambist_a0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_6 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net8939;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_6 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net8939), .TE(1'b0) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net8939), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net8939), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net8939), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net8939), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net8939), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net8939), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net8939), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net8939), .XR(arstz), .Q(rdat[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_6 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_WIDTH5_1 ( clk, arstz, we, wdat, rdat );
  input [4:0] wdat;
  output [4:0] rdat;
  input clk, arstz, we;
  wire   net8957;

  SNPS_CLOCK_GATE_HIGH_glreg_WIDTH5_1 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net8957), .TE(1'b0) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net8957), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net8957), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net8957), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net8957), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net8957), .XR(arstz), .Q(rdat[3]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_WIDTH5_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_WIDTH1_0 ( clk, arstz, we, wdat, rdat );
  input [0:0] wdat;
  output [0:0] rdat;
  input clk, arstz, we;
  wire   n2;

  DFFRQX1 mem_reg_0_ ( .D(n2), .C(clk), .XR(arstz), .Q(rdat[0]) );
  AO22AXL U2 ( .A(we), .B(wdat[0]), .C(rdat[0]), .D(we), .Y(n2) );
endmodule


module regx_a0 ( regx_r, regx_w, di_drposc, di_imposc, di_rd_det, di_stbovp, 
        clk_500k, r_imp_osc, regx_addr, regx_wdat, regx_rdat, regx_hitbst, 
        regx_wrpwm, regx_wrcvc, r_sdischg, r_bistctl, r_bistdat, r_vcomp, 
        r_idacsh, r_cvofsx, r_pwm, regx_wrdac, dac_r_vs, dac_comp, r_dac_en, 
        r_sar_en, r_aopt, r_xtm, r_adummyi, r_bck0, r_bck1, r_i2crout, r_xana, 
        di_xana, lt_gpi, di_tst, bkpt_pc, bkpt_ena, we_twlb, r_vpp_en, 
        r_vpp0v_en, r_otp_pwdn_en, r_otp_wpls, wd_twlb, r_sap, r_twlb, 
        upd_pwrv, ramacc, sse_idle, bus_idle, r_do_ts, r_dpdo_sel, r_dndo_sel, 
        di_ts, detclk, aswclk, atpg_en, di_aswk, clk, rrstz );
  input [6:0] regx_addr;
  input [7:0] regx_wdat;
  output [7:0] regx_rdat;
  output [1:0] regx_hitbst;
  output [1:0] regx_wrpwm;
  output [3:0] regx_wrcvc;
  input [7:0] r_sdischg;
  input [6:0] r_bistctl;
  input [7:0] r_bistdat;
  input [7:0] r_vcomp;
  input [7:0] r_idacsh;
  input [7:0] r_cvofsx;
  input [15:0] r_pwm;
  output [13:0] regx_wrdac;
  input [79:0] dac_r_vs;
  input [9:0] dac_comp;
  input [9:0] r_dac_en;
  input [9:0] r_sar_en;
  output [7:0] r_aopt;
  output [7:0] r_xtm;
  output [7:0] r_adummyi;
  output [7:0] r_bck0;
  output [7:0] r_bck1;
  output [5:0] r_i2crout;
  output [23:0] r_xana;
  input [4:0] di_xana;
  input [3:0] lt_gpi;
  output [14:0] bkpt_pc;
  output [1:0] wd_twlb;
  output [1:0] r_sap;
  input [1:0] r_twlb;
  output [6:0] r_do_ts;
  output [3:0] r_dpdo_sel;
  output [3:0] r_dndo_sel;
  input [4:0] di_aswk;
  input regx_r, regx_w, di_drposc, di_imposc, di_rd_det, di_stbovp, clk_500k,
         di_tst, upd_pwrv, ramacc, sse_idle, bus_idle, di_ts, detclk, aswclk,
         atpg_en, clk, rrstz;
  output r_imp_osc, bkpt_ena, we_twlb, r_vpp_en, r_vpp0v_en, r_otp_pwdn_en,
         r_otp_wpls;
  wire   n109, we_19, we_7, we_5, we_4, reg1F_7, reg1F_6, reg1B_3_, reg10_7_,
         lt_drp, i2c_mode_upd, N8, d_we16, lt_reg1C_0, net8975, n1047, n1048,
         n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
         n1059, n1060, n1061, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n29, n30, n31, n32, n33, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108,
         SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2,
         SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4,
         SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6,
         SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8,
         SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10,
         SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12,
         SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14,
         SYNOPSYS_UNCONNECTED_15, SYNOPSYS_UNCONNECTED_16,
         SYNOPSYS_UNCONNECTED_17, SYNOPSYS_UNCONNECTED_18,
         SYNOPSYS_UNCONNECTED_19, SYNOPSYS_UNCONNECTED_20,
         SYNOPSYS_UNCONNECTED_21, SYNOPSYS_UNCONNECTED_22,
         SYNOPSYS_UNCONNECTED_23, SYNOPSYS_UNCONNECTED_24,
         SYNOPSYS_UNCONNECTED_25, SYNOPSYS_UNCONNECTED_26,
         SYNOPSYS_UNCONNECTED_27, SYNOPSYS_UNCONNECTED_28,
         SYNOPSYS_UNCONNECTED_29, SYNOPSYS_UNCONNECTED_30,
         SYNOPSYS_UNCONNECTED_31, SYNOPSYS_UNCONNECTED_32,
         SYNOPSYS_UNCONNECTED_33, SYNOPSYS_UNCONNECTED_34,
         SYNOPSYS_UNCONNECTED_35, SYNOPSYS_UNCONNECTED_36,
         SYNOPSYS_UNCONNECTED_37, SYNOPSYS_UNCONNECTED_38,
         SYNOPSYS_UNCONNECTED_39, SYNOPSYS_UNCONNECTED_40,
         SYNOPSYS_UNCONNECTED_41, SYNOPSYS_UNCONNECTED_42,
         SYNOPSYS_UNCONNECTED_43, SYNOPSYS_UNCONNECTED_44,
         SYNOPSYS_UNCONNECTED_45, SYNOPSYS_UNCONNECTED_46,
         SYNOPSYS_UNCONNECTED_47, SYNOPSYS_UNCONNECTED_48,
         SYNOPSYS_UNCONNECTED_49, SYNOPSYS_UNCONNECTED_50,
         SYNOPSYS_UNCONNECTED_51, SYNOPSYS_UNCONNECTED_52,
         SYNOPSYS_UNCONNECTED_53, SYNOPSYS_UNCONNECTED_54,
         SYNOPSYS_UNCONNECTED_55, SYNOPSYS_UNCONNECTED_56,
         SYNOPSYS_UNCONNECTED_57, SYNOPSYS_UNCONNECTED_58,
         SYNOPSYS_UNCONNECTED_59, SYNOPSYS_UNCONNECTED_60,
         SYNOPSYS_UNCONNECTED_61, SYNOPSYS_UNCONNECTED_62,
         SYNOPSYS_UNCONNECTED_63, SYNOPSYS_UNCONNECTED_64,
         SYNOPSYS_UNCONNECTED_65, SYNOPSYS_UNCONNECTED_66,
         SYNOPSYS_UNCONNECTED_67, SYNOPSYS_UNCONNECTED_68,
         SYNOPSYS_UNCONNECTED_69, SYNOPSYS_UNCONNECTED_70,
         SYNOPSYS_UNCONNECTED_71, SYNOPSYS_UNCONNECTED_72,
         SYNOPSYS_UNCONNECTED_73, SYNOPSYS_UNCONNECTED_74,
         SYNOPSYS_UNCONNECTED_75, SYNOPSYS_UNCONNECTED_76,
         SYNOPSYS_UNCONNECTED_77, SYNOPSYS_UNCONNECTED_78,
         SYNOPSYS_UNCONNECTED_79, SYNOPSYS_UNCONNECTED_80,
         SYNOPSYS_UNCONNECTED_81, SYNOPSYS_UNCONNECTED_82,
         SYNOPSYS_UNCONNECTED_83, SYNOPSYS_UNCONNECTED_84,
         SYNOPSYS_UNCONNECTED_85, SYNOPSYS_UNCONNECTED_86,
         SYNOPSYS_UNCONNECTED_87, SYNOPSYS_UNCONNECTED_88,
         SYNOPSYS_UNCONNECTED_89, SYNOPSYS_UNCONNECTED_90,
         SYNOPSYS_UNCONNECTED_91, SYNOPSYS_UNCONNECTED_92,
         SYNOPSYS_UNCONNECTED_93, SYNOPSYS_UNCONNECTED_94,
         SYNOPSYS_UNCONNECTED_95, SYNOPSYS_UNCONNECTED_96,
         SYNOPSYS_UNCONNECTED_97, SYNOPSYS_UNCONNECTED_98,
         SYNOPSYS_UNCONNECTED_99, SYNOPSYS_UNCONNECTED_100,
         SYNOPSYS_UNCONNECTED_101, SYNOPSYS_UNCONNECTED_102,
         SYNOPSYS_UNCONNECTED_103, SYNOPSYS_UNCONNECTED_104,
         SYNOPSYS_UNCONNECTED_105, SYNOPSYS_UNCONNECTED_106,
         SYNOPSYS_UNCONNECTED_107, SYNOPSYS_UNCONNECTED_108,
         SYNOPSYS_UNCONNECTED_109, SYNOPSYS_UNCONNECTED_110,
         SYNOPSYS_UNCONNECTED_111, SYNOPSYS_UNCONNECTED_112,
         SYNOPSYS_UNCONNECTED_113, SYNOPSYS_UNCONNECTED_114,
         SYNOPSYS_UNCONNECTED_115, SYNOPSYS_UNCONNECTED_116,
         SYNOPSYS_UNCONNECTED_117, SYNOPSYS_UNCONNECTED_118,
         SYNOPSYS_UNCONNECTED_119, SYNOPSYS_UNCONNECTED_120,
         SYNOPSYS_UNCONNECTED_121, SYNOPSYS_UNCONNECTED_122,
         SYNOPSYS_UNCONNECTED_123, SYNOPSYS_UNCONNECTED_124,
         SYNOPSYS_UNCONNECTED_125, SYNOPSYS_UNCONNECTED_126,
         SYNOPSYS_UNCONNECTED_127, SYNOPSYS_UNCONNECTED_128,
         SYNOPSYS_UNCONNECTED_129, SYNOPSYS_UNCONNECTED_130,
         SYNOPSYS_UNCONNECTED_131, SYNOPSYS_UNCONNECTED_132,
         SYNOPSYS_UNCONNECTED_133, SYNOPSYS_UNCONNECTED_134,
         SYNOPSYS_UNCONNECTED_135, SYNOPSYS_UNCONNECTED_136,
         SYNOPSYS_UNCONNECTED_137, SYNOPSYS_UNCONNECTED_138,
         SYNOPSYS_UNCONNECTED_139, SYNOPSYS_UNCONNECTED_140,
         SYNOPSYS_UNCONNECTED_141, SYNOPSYS_UNCONNECTED_142,
         SYNOPSYS_UNCONNECTED_143, SYNOPSYS_UNCONNECTED_144,
         SYNOPSYS_UNCONNECTED_145, SYNOPSYS_UNCONNECTED_146,
         SYNOPSYS_UNCONNECTED_147, SYNOPSYS_UNCONNECTED_148,
         SYNOPSYS_UNCONNECTED_149, SYNOPSYS_UNCONNECTED_150,
         SYNOPSYS_UNCONNECTED_151, SYNOPSYS_UNCONNECTED_152,
         SYNOPSYS_UNCONNECTED_153, SYNOPSYS_UNCONNECTED_154,
         SYNOPSYS_UNCONNECTED_155, SYNOPSYS_UNCONNECTED_156,
         SYNOPSYS_UNCONNECTED_157, SYNOPSYS_UNCONNECTED_158,
         SYNOPSYS_UNCONNECTED_159, SYNOPSYS_UNCONNECTED_160,
         SYNOPSYS_UNCONNECTED_161, SYNOPSYS_UNCONNECTED_162,
         SYNOPSYS_UNCONNECTED_163, SYNOPSYS_UNCONNECTED_164,
         SYNOPSYS_UNCONNECTED_165, SYNOPSYS_UNCONNECTED_166,
         SYNOPSYS_UNCONNECTED_167, SYNOPSYS_UNCONNECTED_168,
         SYNOPSYS_UNCONNECTED_169, SYNOPSYS_UNCONNECTED_170,
         SYNOPSYS_UNCONNECTED_171, SYNOPSYS_UNCONNECTED_172,
         SYNOPSYS_UNCONNECTED_173, SYNOPSYS_UNCONNECTED_174,
         SYNOPSYS_UNCONNECTED_175, SYNOPSYS_UNCONNECTED_176,
         SYNOPSYS_UNCONNECTED_177, SYNOPSYS_UNCONNECTED_178,
         SYNOPSYS_UNCONNECTED_179, SYNOPSYS_UNCONNECTED_180,
         SYNOPSYS_UNCONNECTED_181, SYNOPSYS_UNCONNECTED_182,
         SYNOPSYS_UNCONNECTED_183, SYNOPSYS_UNCONNECTED_184,
         SYNOPSYS_UNCONNECTED_185, SYNOPSYS_UNCONNECTED_186,
         SYNOPSYS_UNCONNECTED_187, SYNOPSYS_UNCONNECTED_188,
         SYNOPSYS_UNCONNECTED_189, SYNOPSYS_UNCONNECTED_190,
         SYNOPSYS_UNCONNECTED_191, SYNOPSYS_UNCONNECTED_192,
         SYNOPSYS_UNCONNECTED_193, SYNOPSYS_UNCONNECTED_194,
         SYNOPSYS_UNCONNECTED_195, SYNOPSYS_UNCONNECTED_196,
         SYNOPSYS_UNCONNECTED_197, SYNOPSYS_UNCONNECTED_198,
         SYNOPSYS_UNCONNECTED_199, SYNOPSYS_UNCONNECTED_200,
         SYNOPSYS_UNCONNECTED_201, SYNOPSYS_UNCONNECTED_202,
         SYNOPSYS_UNCONNECTED_203, SYNOPSYS_UNCONNECTED_204,
         SYNOPSYS_UNCONNECTED_205, SYNOPSYS_UNCONNECTED_206,
         SYNOPSYS_UNCONNECTED_207, SYNOPSYS_UNCONNECTED_208,
         SYNOPSYS_UNCONNECTED_209, SYNOPSYS_UNCONNECTED_210,
         SYNOPSYS_UNCONNECTED_211, SYNOPSYS_UNCONNECTED_212,
         SYNOPSYS_UNCONNECTED_213, SYNOPSYS_UNCONNECTED_214,
         SYNOPSYS_UNCONNECTED_215, SYNOPSYS_UNCONNECTED_216,
         SYNOPSYS_UNCONNECTED_217, SYNOPSYS_UNCONNECTED_218,
         SYNOPSYS_UNCONNECTED_219, SYNOPSYS_UNCONNECTED_220,
         SYNOPSYS_UNCONNECTED_221, SYNOPSYS_UNCONNECTED_222,
         SYNOPSYS_UNCONNECTED_223, SYNOPSYS_UNCONNECTED_224,
         SYNOPSYS_UNCONNECTED_225, SYNOPSYS_UNCONNECTED_226,
         SYNOPSYS_UNCONNECTED_227, SYNOPSYS_UNCONNECTED_228,
         SYNOPSYS_UNCONNECTED_229, SYNOPSYS_UNCONNECTED_230,
         SYNOPSYS_UNCONNECTED_231, SYNOPSYS_UNCONNECTED_232,
         SYNOPSYS_UNCONNECTED_233, SYNOPSYS_UNCONNECTED_234,
         SYNOPSYS_UNCONNECTED_235, SYNOPSYS_UNCONNECTED_236,
         SYNOPSYS_UNCONNECTED_237, SYNOPSYS_UNCONNECTED_238,
         SYNOPSYS_UNCONNECTED_239, SYNOPSYS_UNCONNECTED_240,
         SYNOPSYS_UNCONNECTED_241, SYNOPSYS_UNCONNECTED_242,
         SYNOPSYS_UNCONNECTED_243, SYNOPSYS_UNCONNECTED_244,
         SYNOPSYS_UNCONNECTED_245, SYNOPSYS_UNCONNECTED_246,
         SYNOPSYS_UNCONNECTED_247, SYNOPSYS_UNCONNECTED_248,
         SYNOPSYS_UNCONNECTED_249, SYNOPSYS_UNCONNECTED_250,
         SYNOPSYS_UNCONNECTED_251, SYNOPSYS_UNCONNECTED_252,
         SYNOPSYS_UNCONNECTED_253, SYNOPSYS_UNCONNECTED_254,
         SYNOPSYS_UNCONNECTED_255, SYNOPSYS_UNCONNECTED_256,
         SYNOPSYS_UNCONNECTED_257, SYNOPSYS_UNCONNECTED_258,
         SYNOPSYS_UNCONNECTED_259, SYNOPSYS_UNCONNECTED_260,
         SYNOPSYS_UNCONNECTED_261, SYNOPSYS_UNCONNECTED_262,
         SYNOPSYS_UNCONNECTED_263, SYNOPSYS_UNCONNECTED_264,
         SYNOPSYS_UNCONNECTED_265, SYNOPSYS_UNCONNECTED_266,
         SYNOPSYS_UNCONNECTED_267, SYNOPSYS_UNCONNECTED_268,
         SYNOPSYS_UNCONNECTED_269, SYNOPSYS_UNCONNECTED_270,
         SYNOPSYS_UNCONNECTED_271, SYNOPSYS_UNCONNECTED_272,
         SYNOPSYS_UNCONNECTED_273, SYNOPSYS_UNCONNECTED_274,
         SYNOPSYS_UNCONNECTED_275, SYNOPSYS_UNCONNECTED_276,
         SYNOPSYS_UNCONNECTED_277, SYNOPSYS_UNCONNECTED_278,
         SYNOPSYS_UNCONNECTED_279, SYNOPSYS_UNCONNECTED_280,
         SYNOPSYS_UNCONNECTED_281, SYNOPSYS_UNCONNECTED_282,
         SYNOPSYS_UNCONNECTED_283, SYNOPSYS_UNCONNECTED_284,
         SYNOPSYS_UNCONNECTED_285, SYNOPSYS_UNCONNECTED_286,
         SYNOPSYS_UNCONNECTED_287, SYNOPSYS_UNCONNECTED_288,
         SYNOPSYS_UNCONNECTED_289, SYNOPSYS_UNCONNECTED_290,
         SYNOPSYS_UNCONNECTED_291, SYNOPSYS_UNCONNECTED_292,
         SYNOPSYS_UNCONNECTED_293, SYNOPSYS_UNCONNECTED_294,
         SYNOPSYS_UNCONNECTED_295, SYNOPSYS_UNCONNECTED_296,
         SYNOPSYS_UNCONNECTED_297, SYNOPSYS_UNCONNECTED_298,
         SYNOPSYS_UNCONNECTED_299, SYNOPSYS_UNCONNECTED_300,
         SYNOPSYS_UNCONNECTED_301, SYNOPSYS_UNCONNECTED_302,
         SYNOPSYS_UNCONNECTED_303, SYNOPSYS_UNCONNECTED_304,
         SYNOPSYS_UNCONNECTED_305, SYNOPSYS_UNCONNECTED_306,
         SYNOPSYS_UNCONNECTED_307, SYNOPSYS_UNCONNECTED_308,
         SYNOPSYS_UNCONNECTED_309, SYNOPSYS_UNCONNECTED_310,
         SYNOPSYS_UNCONNECTED_311, SYNOPSYS_UNCONNECTED_312,
         SYNOPSYS_UNCONNECTED_313, SYNOPSYS_UNCONNECTED_314,
         SYNOPSYS_UNCONNECTED_315, SYNOPSYS_UNCONNECTED_316,
         SYNOPSYS_UNCONNECTED_317, SYNOPSYS_UNCONNECTED_318,
         SYNOPSYS_UNCONNECTED_319, SYNOPSYS_UNCONNECTED_320,
         SYNOPSYS_UNCONNECTED_321, SYNOPSYS_UNCONNECTED_322,
         SYNOPSYS_UNCONNECTED_323, SYNOPSYS_UNCONNECTED_324,
         SYNOPSYS_UNCONNECTED_325, SYNOPSYS_UNCONNECTED_326,
         SYNOPSYS_UNCONNECTED_327, SYNOPSYS_UNCONNECTED_328,
         SYNOPSYS_UNCONNECTED_329, SYNOPSYS_UNCONNECTED_330,
         SYNOPSYS_UNCONNECTED_331, SYNOPSYS_UNCONNECTED_332,
         SYNOPSYS_UNCONNECTED_333, SYNOPSYS_UNCONNECTED_334,
         SYNOPSYS_UNCONNECTED_335, SYNOPSYS_UNCONNECTED_336,
         SYNOPSYS_UNCONNECTED_337, SYNOPSYS_UNCONNECTED_338,
         SYNOPSYS_UNCONNECTED_339, SYNOPSYS_UNCONNECTED_340,
         SYNOPSYS_UNCONNECTED_341, SYNOPSYS_UNCONNECTED_342,
         SYNOPSYS_UNCONNECTED_343, SYNOPSYS_UNCONNECTED_344,
         SYNOPSYS_UNCONNECTED_345, SYNOPSYS_UNCONNECTED_346,
         SYNOPSYS_UNCONNECTED_347, SYNOPSYS_UNCONNECTED_348,
         SYNOPSYS_UNCONNECTED_349, SYNOPSYS_UNCONNECTED_350,
         SYNOPSYS_UNCONNECTED_351, SYNOPSYS_UNCONNECTED_352,
         SYNOPSYS_UNCONNECTED_353, SYNOPSYS_UNCONNECTED_354,
         SYNOPSYS_UNCONNECTED_355, SYNOPSYS_UNCONNECTED_356,
         SYNOPSYS_UNCONNECTED_357, SYNOPSYS_UNCONNECTED_358,
         SYNOPSYS_UNCONNECTED_359, SYNOPSYS_UNCONNECTED_360,
         SYNOPSYS_UNCONNECTED_361, SYNOPSYS_UNCONNECTED_362,
         SYNOPSYS_UNCONNECTED_363, SYNOPSYS_UNCONNECTED_364,
         SYNOPSYS_UNCONNECTED_365, SYNOPSYS_UNCONNECTED_366,
         SYNOPSYS_UNCONNECTED_367, SYNOPSYS_UNCONNECTED_368,
         SYNOPSYS_UNCONNECTED_369, SYNOPSYS_UNCONNECTED_370,
         SYNOPSYS_UNCONNECTED_371, SYNOPSYS_UNCONNECTED_372,
         SYNOPSYS_UNCONNECTED_373, SYNOPSYS_UNCONNECTED_374,
         SYNOPSYS_UNCONNECTED_375, SYNOPSYS_UNCONNECTED_376,
         SYNOPSYS_UNCONNECTED_377, SYNOPSYS_UNCONNECTED_378,
         SYNOPSYS_UNCONNECTED_379, SYNOPSYS_UNCONNECTED_380,
         SYNOPSYS_UNCONNECTED_381, SYNOPSYS_UNCONNECTED_382,
         SYNOPSYS_UNCONNECTED_383, SYNOPSYS_UNCONNECTED_384,
         SYNOPSYS_UNCONNECTED_385, SYNOPSYS_UNCONNECTED_386,
         SYNOPSYS_UNCONNECTED_387, SYNOPSYS_UNCONNECTED_388,
         SYNOPSYS_UNCONNECTED_389, SYNOPSYS_UNCONNECTED_390,
         SYNOPSYS_UNCONNECTED_391, SYNOPSYS_UNCONNECTED_392,
         SYNOPSYS_UNCONNECTED_393, SYNOPSYS_UNCONNECTED_394,
         SYNOPSYS_UNCONNECTED_395, SYNOPSYS_UNCONNECTED_396,
         SYNOPSYS_UNCONNECTED_397, SYNOPSYS_UNCONNECTED_398,
         SYNOPSYS_UNCONNECTED_399, SYNOPSYS_UNCONNECTED_400,
         SYNOPSYS_UNCONNECTED_401, SYNOPSYS_UNCONNECTED_402,
         SYNOPSYS_UNCONNECTED_403, SYNOPSYS_UNCONNECTED_404,
         SYNOPSYS_UNCONNECTED_405, SYNOPSYS_UNCONNECTED_406,
         SYNOPSYS_UNCONNECTED_407, SYNOPSYS_UNCONNECTED_408,
         SYNOPSYS_UNCONNECTED_409, SYNOPSYS_UNCONNECTED_410,
         SYNOPSYS_UNCONNECTED_411, SYNOPSYS_UNCONNECTED_412,
         SYNOPSYS_UNCONNECTED_413, SYNOPSYS_UNCONNECTED_414,
         SYNOPSYS_UNCONNECTED_415, SYNOPSYS_UNCONNECTED_416,
         SYNOPSYS_UNCONNECTED_417, SYNOPSYS_UNCONNECTED_418,
         SYNOPSYS_UNCONNECTED_419, SYNOPSYS_UNCONNECTED_420,
         SYNOPSYS_UNCONNECTED_421, SYNOPSYS_UNCONNECTED_422,
         SYNOPSYS_UNCONNECTED_423, SYNOPSYS_UNCONNECTED_424,
         SYNOPSYS_UNCONNECTED_425, SYNOPSYS_UNCONNECTED_426,
         SYNOPSYS_UNCONNECTED_427, SYNOPSYS_UNCONNECTED_428,
         SYNOPSYS_UNCONNECTED_429, SYNOPSYS_UNCONNECTED_430,
         SYNOPSYS_UNCONNECTED_431, SYNOPSYS_UNCONNECTED_432,
         SYNOPSYS_UNCONNECTED_433, SYNOPSYS_UNCONNECTED_434,
         SYNOPSYS_UNCONNECTED_435, SYNOPSYS_UNCONNECTED_436,
         SYNOPSYS_UNCONNECTED_437, SYNOPSYS_UNCONNECTED_438,
         SYNOPSYS_UNCONNECTED_439, SYNOPSYS_UNCONNECTED_440,
         SYNOPSYS_UNCONNECTED_441, SYNOPSYS_UNCONNECTED_442,
         SYNOPSYS_UNCONNECTED_443, SYNOPSYS_UNCONNECTED_444,
         SYNOPSYS_UNCONNECTED_445, SYNOPSYS_UNCONNECTED_446,
         SYNOPSYS_UNCONNECTED_447, SYNOPSYS_UNCONNECTED_448,
         SYNOPSYS_UNCONNECTED_449, SYNOPSYS_UNCONNECTED_450,
         SYNOPSYS_UNCONNECTED_451, SYNOPSYS_UNCONNECTED_452,
         SYNOPSYS_UNCONNECTED_453, SYNOPSYS_UNCONNECTED_454,
         SYNOPSYS_UNCONNECTED_455, SYNOPSYS_UNCONNECTED_456,
         SYNOPSYS_UNCONNECTED_457, SYNOPSYS_UNCONNECTED_458,
         SYNOPSYS_UNCONNECTED_459, SYNOPSYS_UNCONNECTED_460,
         SYNOPSYS_UNCONNECTED_461, SYNOPSYS_UNCONNECTED_462,
         SYNOPSYS_UNCONNECTED_463, SYNOPSYS_UNCONNECTED_464,
         SYNOPSYS_UNCONNECTED_465, SYNOPSYS_UNCONNECTED_466,
         SYNOPSYS_UNCONNECTED_467, SYNOPSYS_UNCONNECTED_468,
         SYNOPSYS_UNCONNECTED_469, SYNOPSYS_UNCONNECTED_470,
         SYNOPSYS_UNCONNECTED_471, SYNOPSYS_UNCONNECTED_472,
         SYNOPSYS_UNCONNECTED_473, SYNOPSYS_UNCONNECTED_474,
         SYNOPSYS_UNCONNECTED_475, SYNOPSYS_UNCONNECTED_476,
         SYNOPSYS_UNCONNECTED_477, SYNOPSYS_UNCONNECTED_478,
         SYNOPSYS_UNCONNECTED_479, SYNOPSYS_UNCONNECTED_480,
         SYNOPSYS_UNCONNECTED_481, SYNOPSYS_UNCONNECTED_482,
         SYNOPSYS_UNCONNECTED_483, SYNOPSYS_UNCONNECTED_484,
         SYNOPSYS_UNCONNECTED_485, SYNOPSYS_UNCONNECTED_486,
         SYNOPSYS_UNCONNECTED_487, SYNOPSYS_UNCONNECTED_488,
         SYNOPSYS_UNCONNECTED_489, SYNOPSYS_UNCONNECTED_490,
         SYNOPSYS_UNCONNECTED_491, SYNOPSYS_UNCONNECTED_492,
         SYNOPSYS_UNCONNECTED_493, SYNOPSYS_UNCONNECTED_494,
         SYNOPSYS_UNCONNECTED_495, SYNOPSYS_UNCONNECTED_496,
         SYNOPSYS_UNCONNECTED_497, SYNOPSYS_UNCONNECTED_498,
         SYNOPSYS_UNCONNECTED_499, SYNOPSYS_UNCONNECTED_500,
         SYNOPSYS_UNCONNECTED_501, SYNOPSYS_UNCONNECTED_502,
         SYNOPSYS_UNCONNECTED_503, SYNOPSYS_UNCONNECTED_504,
         SYNOPSYS_UNCONNECTED_505, SYNOPSYS_UNCONNECTED_506,
         SYNOPSYS_UNCONNECTED_507, SYNOPSYS_UNCONNECTED_508,
         SYNOPSYS_UNCONNECTED_509, SYNOPSYS_UNCONNECTED_510,
         SYNOPSYS_UNCONNECTED_511, SYNOPSYS_UNCONNECTED_512,
         SYNOPSYS_UNCONNECTED_513, SYNOPSYS_UNCONNECTED_514,
         SYNOPSYS_UNCONNECTED_515, SYNOPSYS_UNCONNECTED_516,
         SYNOPSYS_UNCONNECTED_517, SYNOPSYS_UNCONNECTED_518,
         SYNOPSYS_UNCONNECTED_519, SYNOPSYS_UNCONNECTED_520,
         SYNOPSYS_UNCONNECTED_521, SYNOPSYS_UNCONNECTED_522,
         SYNOPSYS_UNCONNECTED_523, SYNOPSYS_UNCONNECTED_524,
         SYNOPSYS_UNCONNECTED_525, SYNOPSYS_UNCONNECTED_526,
         SYNOPSYS_UNCONNECTED_527, SYNOPSYS_UNCONNECTED_528,
         SYNOPSYS_UNCONNECTED_529, SYNOPSYS_UNCONNECTED_530,
         SYNOPSYS_UNCONNECTED_531, SYNOPSYS_UNCONNECTED_532,
         SYNOPSYS_UNCONNECTED_533, SYNOPSYS_UNCONNECTED_534,
         SYNOPSYS_UNCONNECTED_535, SYNOPSYS_UNCONNECTED_536,
         SYNOPSYS_UNCONNECTED_537, SYNOPSYS_UNCONNECTED_538,
         SYNOPSYS_UNCONNECTED_539, SYNOPSYS_UNCONNECTED_540,
         SYNOPSYS_UNCONNECTED_541, SYNOPSYS_UNCONNECTED_542,
         SYNOPSYS_UNCONNECTED_543, SYNOPSYS_UNCONNECTED_544,
         SYNOPSYS_UNCONNECTED_545, SYNOPSYS_UNCONNECTED_546,
         SYNOPSYS_UNCONNECTED_547, SYNOPSYS_UNCONNECTED_548,
         SYNOPSYS_UNCONNECTED_549, SYNOPSYS_UNCONNECTED_550,
         SYNOPSYS_UNCONNECTED_551, SYNOPSYS_UNCONNECTED_552,
         SYNOPSYS_UNCONNECTED_553, SYNOPSYS_UNCONNECTED_554,
         SYNOPSYS_UNCONNECTED_555, SYNOPSYS_UNCONNECTED_556,
         SYNOPSYS_UNCONNECTED_557, SYNOPSYS_UNCONNECTED_558,
         SYNOPSYS_UNCONNECTED_559, SYNOPSYS_UNCONNECTED_560,
         SYNOPSYS_UNCONNECTED_561, SYNOPSYS_UNCONNECTED_562,
         SYNOPSYS_UNCONNECTED_563, SYNOPSYS_UNCONNECTED_564,
         SYNOPSYS_UNCONNECTED_565, SYNOPSYS_UNCONNECTED_566,
         SYNOPSYS_UNCONNECTED_567, SYNOPSYS_UNCONNECTED_568,
         SYNOPSYS_UNCONNECTED_569, SYNOPSYS_UNCONNECTED_570,
         SYNOPSYS_UNCONNECTED_571, SYNOPSYS_UNCONNECTED_572,
         SYNOPSYS_UNCONNECTED_573, SYNOPSYS_UNCONNECTED_574,
         SYNOPSYS_UNCONNECTED_575, SYNOPSYS_UNCONNECTED_576,
         SYNOPSYS_UNCONNECTED_577, SYNOPSYS_UNCONNECTED_578,
         SYNOPSYS_UNCONNECTED_579, SYNOPSYS_UNCONNECTED_580,
         SYNOPSYS_UNCONNECTED_581, SYNOPSYS_UNCONNECTED_582,
         SYNOPSYS_UNCONNECTED_583, SYNOPSYS_UNCONNECTED_584,
         SYNOPSYS_UNCONNECTED_585, SYNOPSYS_UNCONNECTED_586,
         SYNOPSYS_UNCONNECTED_587, SYNOPSYS_UNCONNECTED_588,
         SYNOPSYS_UNCONNECTED_589, SYNOPSYS_UNCONNECTED_590,
         SYNOPSYS_UNCONNECTED_591, SYNOPSYS_UNCONNECTED_592,
         SYNOPSYS_UNCONNECTED_593, SYNOPSYS_UNCONNECTED_594,
         SYNOPSYS_UNCONNECTED_595, SYNOPSYS_UNCONNECTED_596,
         SYNOPSYS_UNCONNECTED_597, SYNOPSYS_UNCONNECTED_598,
         SYNOPSYS_UNCONNECTED_599, SYNOPSYS_UNCONNECTED_600,
         SYNOPSYS_UNCONNECTED_601, SYNOPSYS_UNCONNECTED_602,
         SYNOPSYS_UNCONNECTED_603, SYNOPSYS_UNCONNECTED_604,
         SYNOPSYS_UNCONNECTED_605, SYNOPSYS_UNCONNECTED_606,
         SYNOPSYS_UNCONNECTED_607, SYNOPSYS_UNCONNECTED_608,
         SYNOPSYS_UNCONNECTED_609, SYNOPSYS_UNCONNECTED_610,
         SYNOPSYS_UNCONNECTED_611, SYNOPSYS_UNCONNECTED_612,
         SYNOPSYS_UNCONNECTED_613, SYNOPSYS_UNCONNECTED_614,
         SYNOPSYS_UNCONNECTED_615, SYNOPSYS_UNCONNECTED_616,
         SYNOPSYS_UNCONNECTED_617, SYNOPSYS_UNCONNECTED_618,
         SYNOPSYS_UNCONNECTED_619, SYNOPSYS_UNCONNECTED_620,
         SYNOPSYS_UNCONNECTED_621, SYNOPSYS_UNCONNECTED_622,
         SYNOPSYS_UNCONNECTED_623, SYNOPSYS_UNCONNECTED_624,
         SYNOPSYS_UNCONNECTED_625, SYNOPSYS_UNCONNECTED_626,
         SYNOPSYS_UNCONNECTED_627, SYNOPSYS_UNCONNECTED_628,
         SYNOPSYS_UNCONNECTED_629, SYNOPSYS_UNCONNECTED_630,
         SYNOPSYS_UNCONNECTED_631, SYNOPSYS_UNCONNECTED_632,
         SYNOPSYS_UNCONNECTED_633, SYNOPSYS_UNCONNECTED_634,
         SYNOPSYS_UNCONNECTED_635, SYNOPSYS_UNCONNECTED_636,
         SYNOPSYS_UNCONNECTED_637, SYNOPSYS_UNCONNECTED_638,
         SYNOPSYS_UNCONNECTED_639, SYNOPSYS_UNCONNECTED_640,
         SYNOPSYS_UNCONNECTED_641, SYNOPSYS_UNCONNECTED_642,
         SYNOPSYS_UNCONNECTED_643, SYNOPSYS_UNCONNECTED_644,
         SYNOPSYS_UNCONNECTED_645, SYNOPSYS_UNCONNECTED_646,
         SYNOPSYS_UNCONNECTED_647, SYNOPSYS_UNCONNECTED_648,
         SYNOPSYS_UNCONNECTED_649, SYNOPSYS_UNCONNECTED_650,
         SYNOPSYS_UNCONNECTED_651, SYNOPSYS_UNCONNECTED_652,
         SYNOPSYS_UNCONNECTED_653, SYNOPSYS_UNCONNECTED_654,
         SYNOPSYS_UNCONNECTED_655, SYNOPSYS_UNCONNECTED_656,
         SYNOPSYS_UNCONNECTED_657, SYNOPSYS_UNCONNECTED_658,
         SYNOPSYS_UNCONNECTED_659, SYNOPSYS_UNCONNECTED_660,
         SYNOPSYS_UNCONNECTED_661, SYNOPSYS_UNCONNECTED_662,
         SYNOPSYS_UNCONNECTED_663, SYNOPSYS_UNCONNECTED_664,
         SYNOPSYS_UNCONNECTED_665, SYNOPSYS_UNCONNECTED_666,
         SYNOPSYS_UNCONNECTED_667, SYNOPSYS_UNCONNECTED_668,
         SYNOPSYS_UNCONNECTED_669, SYNOPSYS_UNCONNECTED_670,
         SYNOPSYS_UNCONNECTED_671, SYNOPSYS_UNCONNECTED_672,
         SYNOPSYS_UNCONNECTED_673, SYNOPSYS_UNCONNECTED_674,
         SYNOPSYS_UNCONNECTED_675, SYNOPSYS_UNCONNECTED_676,
         SYNOPSYS_UNCONNECTED_677, SYNOPSYS_UNCONNECTED_678,
         SYNOPSYS_UNCONNECTED_679, SYNOPSYS_UNCONNECTED_680,
         SYNOPSYS_UNCONNECTED_681, SYNOPSYS_UNCONNECTED_682,
         SYNOPSYS_UNCONNECTED_683, SYNOPSYS_UNCONNECTED_684,
         SYNOPSYS_UNCONNECTED_685, SYNOPSYS_UNCONNECTED_686,
         SYNOPSYS_UNCONNECTED_687, SYNOPSYS_UNCONNECTED_688,
         SYNOPSYS_UNCONNECTED_689, SYNOPSYS_UNCONNECTED_690,
         SYNOPSYS_UNCONNECTED_691, SYNOPSYS_UNCONNECTED_692,
         SYNOPSYS_UNCONNECTED_693, SYNOPSYS_UNCONNECTED_694,
         SYNOPSYS_UNCONNECTED_695, SYNOPSYS_UNCONNECTED_696,
         SYNOPSYS_UNCONNECTED_697, SYNOPSYS_UNCONNECTED_698,
         SYNOPSYS_UNCONNECTED_699, SYNOPSYS_UNCONNECTED_700,
         SYNOPSYS_UNCONNECTED_701, SYNOPSYS_UNCONNECTED_702,
         SYNOPSYS_UNCONNECTED_703, SYNOPSYS_UNCONNECTED_704,
         SYNOPSYS_UNCONNECTED_705, SYNOPSYS_UNCONNECTED_706,
         SYNOPSYS_UNCONNECTED_707, SYNOPSYS_UNCONNECTED_708,
         SYNOPSYS_UNCONNECTED_709, SYNOPSYS_UNCONNECTED_710,
         SYNOPSYS_UNCONNECTED_711, SYNOPSYS_UNCONNECTED_712,
         SYNOPSYS_UNCONNECTED_713, SYNOPSYS_UNCONNECTED_714,
         SYNOPSYS_UNCONNECTED_715, SYNOPSYS_UNCONNECTED_716,
         SYNOPSYS_UNCONNECTED_717, SYNOPSYS_UNCONNECTED_718,
         SYNOPSYS_UNCONNECTED_719, SYNOPSYS_UNCONNECTED_720,
         SYNOPSYS_UNCONNECTED_721, SYNOPSYS_UNCONNECTED_722,
         SYNOPSYS_UNCONNECTED_723, SYNOPSYS_UNCONNECTED_724,
         SYNOPSYS_UNCONNECTED_725, SYNOPSYS_UNCONNECTED_726,
         SYNOPSYS_UNCONNECTED_727, SYNOPSYS_UNCONNECTED_728,
         SYNOPSYS_UNCONNECTED_729, SYNOPSYS_UNCONNECTED_730,
         SYNOPSYS_UNCONNECTED_731, SYNOPSYS_UNCONNECTED_732,
         SYNOPSYS_UNCONNECTED_733, SYNOPSYS_UNCONNECTED_734,
         SYNOPSYS_UNCONNECTED_735, SYNOPSYS_UNCONNECTED_736,
         SYNOPSYS_UNCONNECTED_737, SYNOPSYS_UNCONNECTED_738,
         SYNOPSYS_UNCONNECTED_739, SYNOPSYS_UNCONNECTED_740,
         SYNOPSYS_UNCONNECTED_741, SYNOPSYS_UNCONNECTED_742,
         SYNOPSYS_UNCONNECTED_743, SYNOPSYS_UNCONNECTED_744,
         SYNOPSYS_UNCONNECTED_745, SYNOPSYS_UNCONNECTED_746,
         SYNOPSYS_UNCONNECTED_747, SYNOPSYS_UNCONNECTED_748,
         SYNOPSYS_UNCONNECTED_749, SYNOPSYS_UNCONNECTED_750,
         SYNOPSYS_UNCONNECTED_751, SYNOPSYS_UNCONNECTED_752,
         SYNOPSYS_UNCONNECTED_753, SYNOPSYS_UNCONNECTED_754,
         SYNOPSYS_UNCONNECTED_755, SYNOPSYS_UNCONNECTED_756,
         SYNOPSYS_UNCONNECTED_757, SYNOPSYS_UNCONNECTED_758,
         SYNOPSYS_UNCONNECTED_759, SYNOPSYS_UNCONNECTED_760,
         SYNOPSYS_UNCONNECTED_761, SYNOPSYS_UNCONNECTED_762,
         SYNOPSYS_UNCONNECTED_763, SYNOPSYS_UNCONNECTED_764,
         SYNOPSYS_UNCONNECTED_765, SYNOPSYS_UNCONNECTED_766,
         SYNOPSYS_UNCONNECTED_767, SYNOPSYS_UNCONNECTED_768,
         SYNOPSYS_UNCONNECTED_769, SYNOPSYS_UNCONNECTED_770,
         SYNOPSYS_UNCONNECTED_771, SYNOPSYS_UNCONNECTED_772,
         SYNOPSYS_UNCONNECTED_773, SYNOPSYS_UNCONNECTED_774,
         SYNOPSYS_UNCONNECTED_775, SYNOPSYS_UNCONNECTED_776,
         SYNOPSYS_UNCONNECTED_777, SYNOPSYS_UNCONNECTED_778,
         SYNOPSYS_UNCONNECTED_779, SYNOPSYS_UNCONNECTED_780,
         SYNOPSYS_UNCONNECTED_781, SYNOPSYS_UNCONNECTED_782,
         SYNOPSYS_UNCONNECTED_783, SYNOPSYS_UNCONNECTED_784,
         SYNOPSYS_UNCONNECTED_785, SYNOPSYS_UNCONNECTED_786,
         SYNOPSYS_UNCONNECTED_787, SYNOPSYS_UNCONNECTED_788,
         SYNOPSYS_UNCONNECTED_789, SYNOPSYS_UNCONNECTED_790,
         SYNOPSYS_UNCONNECTED_791, SYNOPSYS_UNCONNECTED_792,
         SYNOPSYS_UNCONNECTED_793, SYNOPSYS_UNCONNECTED_794,
         SYNOPSYS_UNCONNECTED_795, SYNOPSYS_UNCONNECTED_796,
         SYNOPSYS_UNCONNECTED_797, SYNOPSYS_UNCONNECTED_798,
         SYNOPSYS_UNCONNECTED_799, SYNOPSYS_UNCONNECTED_800,
         SYNOPSYS_UNCONNECTED_801, SYNOPSYS_UNCONNECTED_802,
         SYNOPSYS_UNCONNECTED_803, SYNOPSYS_UNCONNECTED_804,
         SYNOPSYS_UNCONNECTED_805, SYNOPSYS_UNCONNECTED_806,
         SYNOPSYS_UNCONNECTED_807, SYNOPSYS_UNCONNECTED_808,
         SYNOPSYS_UNCONNECTED_809, SYNOPSYS_UNCONNECTED_810,
         SYNOPSYS_UNCONNECTED_811, SYNOPSYS_UNCONNECTED_812,
         SYNOPSYS_UNCONNECTED_813, SYNOPSYS_UNCONNECTED_814,
         SYNOPSYS_UNCONNECTED_815, SYNOPSYS_UNCONNECTED_816,
         SYNOPSYS_UNCONNECTED_817, SYNOPSYS_UNCONNECTED_818,
         SYNOPSYS_UNCONNECTED_819, SYNOPSYS_UNCONNECTED_820,
         SYNOPSYS_UNCONNECTED_821, SYNOPSYS_UNCONNECTED_822,
         SYNOPSYS_UNCONNECTED_823, SYNOPSYS_UNCONNECTED_824,
         SYNOPSYS_UNCONNECTED_825, SYNOPSYS_UNCONNECTED_826,
         SYNOPSYS_UNCONNECTED_827, SYNOPSYS_UNCONNECTED_828,
         SYNOPSYS_UNCONNECTED_829, SYNOPSYS_UNCONNECTED_830,
         SYNOPSYS_UNCONNECTED_831, SYNOPSYS_UNCONNECTED_832,
         SYNOPSYS_UNCONNECTED_833, SYNOPSYS_UNCONNECTED_834,
         SYNOPSYS_UNCONNECTED_835, SYNOPSYS_UNCONNECTED_836,
         SYNOPSYS_UNCONNECTED_837, SYNOPSYS_UNCONNECTED_838,
         SYNOPSYS_UNCONNECTED_839, SYNOPSYS_UNCONNECTED_840,
         SYNOPSYS_UNCONNECTED_841, SYNOPSYS_UNCONNECTED_842,
         SYNOPSYS_UNCONNECTED_843, SYNOPSYS_UNCONNECTED_844,
         SYNOPSYS_UNCONNECTED_845, SYNOPSYS_UNCONNECTED_846,
         SYNOPSYS_UNCONNECTED_847, SYNOPSYS_UNCONNECTED_848,
         SYNOPSYS_UNCONNECTED_849, SYNOPSYS_UNCONNECTED_850,
         SYNOPSYS_UNCONNECTED_851, SYNOPSYS_UNCONNECTED_852,
         SYNOPSYS_UNCONNECTED_853, SYNOPSYS_UNCONNECTED_854,
         SYNOPSYS_UNCONNECTED_855, SYNOPSYS_UNCONNECTED_856,
         SYNOPSYS_UNCONNECTED_857, SYNOPSYS_UNCONNECTED_858,
         SYNOPSYS_UNCONNECTED_859, SYNOPSYS_UNCONNECTED_860,
         SYNOPSYS_UNCONNECTED_861, SYNOPSYS_UNCONNECTED_862,
         SYNOPSYS_UNCONNECTED_863, SYNOPSYS_UNCONNECTED_864,
         SYNOPSYS_UNCONNECTED_865, SYNOPSYS_UNCONNECTED_866,
         SYNOPSYS_UNCONNECTED_867, SYNOPSYS_UNCONNECTED_868,
         SYNOPSYS_UNCONNECTED_869, SYNOPSYS_UNCONNECTED_870,
         SYNOPSYS_UNCONNECTED_871, SYNOPSYS_UNCONNECTED_872,
         SYNOPSYS_UNCONNECTED_873, SYNOPSYS_UNCONNECTED_874,
         SYNOPSYS_UNCONNECTED_875, SYNOPSYS_UNCONNECTED_876,
         SYNOPSYS_UNCONNECTED_877, SYNOPSYS_UNCONNECTED_878,
         SYNOPSYS_UNCONNECTED_879, SYNOPSYS_UNCONNECTED_880,
         SYNOPSYS_UNCONNECTED_881, SYNOPSYS_UNCONNECTED_882,
         SYNOPSYS_UNCONNECTED_883, SYNOPSYS_UNCONNECTED_884,
         SYNOPSYS_UNCONNECTED_885, SYNOPSYS_UNCONNECTED_886,
         SYNOPSYS_UNCONNECTED_887, SYNOPSYS_UNCONNECTED_888,
         SYNOPSYS_UNCONNECTED_889, SYNOPSYS_UNCONNECTED_890,
         SYNOPSYS_UNCONNECTED_891, SYNOPSYS_UNCONNECTED_892,
         SYNOPSYS_UNCONNECTED_893, SYNOPSYS_UNCONNECTED_894,
         SYNOPSYS_UNCONNECTED_895, SYNOPSYS_UNCONNECTED_896,
         SYNOPSYS_UNCONNECTED_897, SYNOPSYS_UNCONNECTED_898,
         SYNOPSYS_UNCONNECTED_899, SYNOPSYS_UNCONNECTED_900,
         SYNOPSYS_UNCONNECTED_901, SYNOPSYS_UNCONNECTED_902,
         SYNOPSYS_UNCONNECTED_903, SYNOPSYS_UNCONNECTED_904,
         SYNOPSYS_UNCONNECTED_905, SYNOPSYS_UNCONNECTED_906,
         SYNOPSYS_UNCONNECTED_907, SYNOPSYS_UNCONNECTED_908,
         SYNOPSYS_UNCONNECTED_909, SYNOPSYS_UNCONNECTED_910,
         SYNOPSYS_UNCONNECTED_911, SYNOPSYS_UNCONNECTED_912,
         SYNOPSYS_UNCONNECTED_913, SYNOPSYS_UNCONNECTED_914,
         SYNOPSYS_UNCONNECTED_915, SYNOPSYS_UNCONNECTED_916,
         SYNOPSYS_UNCONNECTED_917, SYNOPSYS_UNCONNECTED_918,
         SYNOPSYS_UNCONNECTED_919, SYNOPSYS_UNCONNECTED_920,
         SYNOPSYS_UNCONNECTED_921, SYNOPSYS_UNCONNECTED_922,
         SYNOPSYS_UNCONNECTED_923, SYNOPSYS_UNCONNECTED_924,
         SYNOPSYS_UNCONNECTED_925, SYNOPSYS_UNCONNECTED_926,
         SYNOPSYS_UNCONNECTED_927, SYNOPSYS_UNCONNECTED_928,
         SYNOPSYS_UNCONNECTED_929, SYNOPSYS_UNCONNECTED_930,
         SYNOPSYS_UNCONNECTED_931, SYNOPSYS_UNCONNECTED_932,
         SYNOPSYS_UNCONNECTED_933, SYNOPSYS_UNCONNECTED_934,
         SYNOPSYS_UNCONNECTED_935, SYNOPSYS_UNCONNECTED_936,
         SYNOPSYS_UNCONNECTED_937, SYNOPSYS_UNCONNECTED_938,
         SYNOPSYS_UNCONNECTED_939, SYNOPSYS_UNCONNECTED_940,
         SYNOPSYS_UNCONNECTED_941, SYNOPSYS_UNCONNECTED_942,
         SYNOPSYS_UNCONNECTED_943, SYNOPSYS_UNCONNECTED_944,
         SYNOPSYS_UNCONNECTED_945, SYNOPSYS_UNCONNECTED_946,
         SYNOPSYS_UNCONNECTED_947, SYNOPSYS_UNCONNECTED_948,
         SYNOPSYS_UNCONNECTED_949, SYNOPSYS_UNCONNECTED_950,
         SYNOPSYS_UNCONNECTED_951, SYNOPSYS_UNCONNECTED_952,
         SYNOPSYS_UNCONNECTED_953, SYNOPSYS_UNCONNECTED_954,
         SYNOPSYS_UNCONNECTED_955, SYNOPSYS_UNCONNECTED_956,
         SYNOPSYS_UNCONNECTED_957, SYNOPSYS_UNCONNECTED_958,
         SYNOPSYS_UNCONNECTED_959, SYNOPSYS_UNCONNECTED_960,
         SYNOPSYS_UNCONNECTED_961, SYNOPSYS_UNCONNECTED_962,
         SYNOPSYS_UNCONNECTED_963, SYNOPSYS_UNCONNECTED_964,
         SYNOPSYS_UNCONNECTED_965, SYNOPSYS_UNCONNECTED_966,
         SYNOPSYS_UNCONNECTED_967, SYNOPSYS_UNCONNECTED_968,
         SYNOPSYS_UNCONNECTED_969, SYNOPSYS_UNCONNECTED_970,
         SYNOPSYS_UNCONNECTED_971, SYNOPSYS_UNCONNECTED_972,
         SYNOPSYS_UNCONNECTED_973, SYNOPSYS_UNCONNECTED_974,
         SYNOPSYS_UNCONNECTED_975, SYNOPSYS_UNCONNECTED_976,
         SYNOPSYS_UNCONNECTED_977, SYNOPSYS_UNCONNECTED_978,
         SYNOPSYS_UNCONNECTED_979, SYNOPSYS_UNCONNECTED_980,
         SYNOPSYS_UNCONNECTED_981, SYNOPSYS_UNCONNECTED_982,
         SYNOPSYS_UNCONNECTED_983, SYNOPSYS_UNCONNECTED_984,
         SYNOPSYS_UNCONNECTED_985, SYNOPSYS_UNCONNECTED_986,
         SYNOPSYS_UNCONNECTED_987, SYNOPSYS_UNCONNECTED_988,
         SYNOPSYS_UNCONNECTED_989, SYNOPSYS_UNCONNECTED_990,
         SYNOPSYS_UNCONNECTED_991, SYNOPSYS_UNCONNECTED_992,
         SYNOPSYS_UNCONNECTED_993, SYNOPSYS_UNCONNECTED_994,
         SYNOPSYS_UNCONNECTED_995, SYNOPSYS_UNCONNECTED_996,
         SYNOPSYS_UNCONNECTED_997, SYNOPSYS_UNCONNECTED_998,
         SYNOPSYS_UNCONNECTED_999, SYNOPSYS_UNCONNECTED_1000,
         SYNOPSYS_UNCONNECTED_1001, SYNOPSYS_UNCONNECTED_1002,
         SYNOPSYS_UNCONNECTED_1003, SYNOPSYS_UNCONNECTED_1004,
         SYNOPSYS_UNCONNECTED_1005, SYNOPSYS_UNCONNECTED_1006,
         SYNOPSYS_UNCONNECTED_1007, SYNOPSYS_UNCONNECTED_1008,
         SYNOPSYS_UNCONNECTED_1009, SYNOPSYS_UNCONNECTED_1010,
         SYNOPSYS_UNCONNECTED_1011, SYNOPSYS_UNCONNECTED_1012,
         SYNOPSYS_UNCONNECTED_1013, SYNOPSYS_UNCONNECTED_1014,
         SYNOPSYS_UNCONNECTED_1015, SYNOPSYS_UNCONNECTED_1016;
  wire   [30:23] we;
  wire   [6:0] d_regx_addr;
  wire   [4:0] reg1F;
  wire   [3:2] reg1E;
  wire   [3:0] reg14;
  wire   [3:0] d_lt_gpi;
  wire   [5:0] lt_reg15_5_0;
  wire   [5:0] i2c_mode_wdat;
  wire   [5:0] d_lt_aswk;
  wire   [5:0] lt_aswk;
  wire   [7:0] wd18;

  glreg_a0_18 u0_reg04 ( .clk(clk), .arstz(n38), .we(we_4), .wdat({n18, n8, 
        n16, n13, n5, n22, n10, n24}), .rdat(r_bck0) );
  glreg_a0_17 u0_reg05 ( .clk(clk), .arstz(n39), .we(we_5), .wdat({n19, n8, 
        n15, n12, n4, n22, n10, n24}), .rdat(r_bck1) );
  glreg_a0_16 u0_reg07 ( .clk(clk), .arstz(n40), .we(we_7), .wdat({n18, n7, 
        n15, n12, n5, regx_wdat[2], wd_twlb[1], n24}), .rdat(r_adummyi) );
  glreg_WIDTH1_2 u0_reg10 ( .clk(clk), .arstz(n42), .we(1'b1), .wdat(ramacc), 
        .rdat(reg10_7_) );
  glreg_6_00000002 u0_reg12 ( .clk(clk), .arstz(n51), .we(we_twlb), .wdat({n19, 
        n8, n16, n13, n5, n21}), .rdat({r_vpp_en, r_vpp0v_en, r_otp_pwdn_en, 
        r_otp_wpls, r_sap}) );
  glreg_a0_15 u0_reg13 ( .clk(clk), .arstz(n41), .we(we_19), .wdat({n19, n8, 
        n16, n13, n5, n22, n10, wd_twlb[0]}), .rdat({r_dpdo_sel, r_dndo_sel})
         );
  glreg_WIDTH6_1 u0_reg15 ( .clk(clk), .arstz(n55), .we(n25), .wdat({n16, n13, 
        n5, n22, n10, wd_twlb[0]}), .rdat(lt_reg15_5_0) );
  glreg_WIDTH6_0 u1_reg15 ( .clk(clk), .arstz(n54), .we(i2c_mode_upd), .wdat(
        i2c_mode_wdat), .rdat({n109, r_i2crout[4:0]}) );
  glreg_a0_14 u0_reg17 ( .clk(clk), .arstz(n42), .we(we[23]), .wdat({n19, n7, 
        n15, n12, n4, n21, n10, n24}), .rdat(r_aopt) );
  glreg_a0_13 u0_tmp18 ( .clk(clk), .arstz(n43), .we(we[24]), .wdat({n18, n7, 
        n16, n13, n5, n21, regx_wdat[1], n24}), .rdat(wd18) );
  glreg_a0_12 u0_reg18 ( .clk(clk), .arstz(n44), .we(we[25]), .wdat(wd18), 
        .rdat(bkpt_pc[7:0]) );
  glreg_a0_11 u0_reg19 ( .clk(clk), .arstz(n45), .we(we[25]), .wdat({n19, n8, 
        n16, n13, n5, n22, wd_twlb[1], regx_wdat[0]}), .rdat({bkpt_ena, 
        bkpt_pc[14:8]}) );
  glreg_a0_10 u0_reg1A ( .clk(clk), .arstz(n46), .we(we[26]), .wdat({n19, n8, 
        n16, n13, n5, n22, n10, wd_twlb[0]}), .rdat(r_xtm) );
  dbnc_WIDTH2_TIMEOUT2_7 u0_ts_db ( .o_dbc(reg1B_3_), .o_chg(), .i_org(di_ts), 
        .clk(clk), .rstz(n57) );
  glreg_WIDTH7_0 u0_reg1B ( .clk(clk), .arstz(n50), .we(we[27]), .wdat({n19, 
        n8, n15, n12, n22, n10, n24}), .rdat(r_do_ts) );
  glreg_WIDTH1_1 u1_reg1C ( .clk(clk), .arstz(n38), .we(upd_pwrv), .wdat(
        lt_reg1C_0), .rdat(r_xana[0]) );
  glreg_a0_9 u0_reg1C ( .clk(clk), .arstz(n49), .we(we[28]), .wdat({n18, n7, 
        n16, n13, n4, n21, regx_wdat[1], n24}), .rdat({r_xana[7:1], lt_reg1C_0}) );
  glreg_a0_8 u0_reg1D ( .clk(clk), .arstz(n47), .we(we[29]), .wdat({n19, n8, 
        n16, n13, n5, n22, wd_twlb}), .rdat(r_xana[15:8]) );
  glreg_a0_7 u0_reg1E ( .clk(clk), .arstz(n48), .we(we[30]), .wdat({n19, n8, 
        n16, n13, n5, n22, n10, wd_twlb[0]}), .rdat({r_xana[23], r_imp_osc, 
        r_xana[21:20], reg1E, r_xana[17:16]}) );
  dbnc_WIDTH2_TIMEOUT2_6 u0_dosc_db ( .o_dbc(reg14[1]), .o_chg(), .i_org(
        di_imposc), .clk(clk), .rstz(n54) );
  dbnc_WIDTH2_TIMEOUT2_5 u0_iosc_db ( .o_dbc(reg14[2]), .o_chg(), .i_org(
        di_drposc), .clk(clk), .rstz(n56) );
  dbnc_WIDTH2_TIMEOUT2_4 u0_xana_db ( .o_dbc(reg1F[0]), .o_chg(), .i_org(
        di_xana[0]), .clk(clk), .rstz(n57) );
  dbnc_WIDTH2_TIMEOUT2_3 u1_xana_db ( .o_dbc(reg1F[1]), .o_chg(), .i_org(
        di_xana[1]), .clk(clk), .rstz(rrstz) );
  dbnc_WIDTH2_TIMEOUT2_2 u2_xana_db ( .o_dbc(reg1F[2]), .o_chg(), .i_org(
        di_xana[2]), .clk(clk), .rstz(n55) );
  dbnc_WIDTH2_TIMEOUT2_1 u3_xana_db ( .o_dbc(reg1F[3]), .o_chg(), .i_org(
        di_xana[3]), .clk(clk), .rstz(n56) );
  dbnc_WIDTH2_TIMEOUT2_0 u4_xana_db ( .o_dbc(reg1F[4]), .o_chg(), .i_org(
        di_xana[4]), .clk(clk), .rstz(n51) );
  dbnc_a0_1 u0_sbov_db ( .o_dbc(reg1F_6), .o_chg(), .i_org(di_stbovp), .clk(
        clk_500k), .rstz(n52) );
  dbnc_a0_0 u0_rdet_db ( .o_dbc(reg1F_7), .o_chg(), .i_org(di_rd_det), .clk(
        clk_500k), .rstz(n53) );
  SNPS_CLOCK_GATE_HIGH_regx_a0 clk_gate_d_lt_gpi_reg ( .CLK(clk), .EN(n60), 
        .ENCLK(net8975), .TE(1'b0) );
  regx_a0_DW_rightsh_0 srl_66 ( .A({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        dac_comp[9:8], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, r_sar_en[9:8], 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, r_dac_en[9:8], 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        dac_comp[7:0], r_sar_en[7:0], r_dac_en[7:0], dac_r_vs[63:0], 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        dac_r_vs[79:64], reg1F_7, reg1F_6, 1'b0, reg1F, r_xana[23], r_imp_osc, 
        r_xana[21:20], reg1E, r_xana[17:0], r_do_ts[6:3], reg1B_3_, 
        r_do_ts[2:0], r_xtm, bkpt_ena, bkpt_pc, r_aopt, 1'b0, 1'b0, d_lt_aswk, 
        sse_idle, 1'b0, r_i2crout, d_lt_gpi, reg14, r_dpdo_sel, r_dndo_sel, 
        r_vpp_en, r_vpp0v_en, r_otp_pwdn_en, r_otp_wpls, r_sap, r_twlb, 
        r_bistdat, reg10_7_, r_bistctl, r_sdischg, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        r_pwm, r_adummyi, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        r_bck1, r_bck0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        r_cvofsx, r_idacsh, r_vcomp}), .DATA_TC(1'b0), .SH({d_regx_addr, 1'b0, 
        1'b0, 1'b0}), .B({SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2, 
        SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5, 
        SYNOPSYS_UNCONNECTED_6, SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8, 
        SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10, 
        SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12, 
        SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14, 
        SYNOPSYS_UNCONNECTED_15, SYNOPSYS_UNCONNECTED_16, 
        SYNOPSYS_UNCONNECTED_17, SYNOPSYS_UNCONNECTED_18, 
        SYNOPSYS_UNCONNECTED_19, SYNOPSYS_UNCONNECTED_20, 
        SYNOPSYS_UNCONNECTED_21, SYNOPSYS_UNCONNECTED_22, 
        SYNOPSYS_UNCONNECTED_23, SYNOPSYS_UNCONNECTED_24, 
        SYNOPSYS_UNCONNECTED_25, SYNOPSYS_UNCONNECTED_26, 
        SYNOPSYS_UNCONNECTED_27, SYNOPSYS_UNCONNECTED_28, 
        SYNOPSYS_UNCONNECTED_29, SYNOPSYS_UNCONNECTED_30, 
        SYNOPSYS_UNCONNECTED_31, SYNOPSYS_UNCONNECTED_32, 
        SYNOPSYS_UNCONNECTED_33, SYNOPSYS_UNCONNECTED_34, 
        SYNOPSYS_UNCONNECTED_35, SYNOPSYS_UNCONNECTED_36, 
        SYNOPSYS_UNCONNECTED_37, SYNOPSYS_UNCONNECTED_38, 
        SYNOPSYS_UNCONNECTED_39, SYNOPSYS_UNCONNECTED_40, 
        SYNOPSYS_UNCONNECTED_41, SYNOPSYS_UNCONNECTED_42, 
        SYNOPSYS_UNCONNECTED_43, SYNOPSYS_UNCONNECTED_44, 
        SYNOPSYS_UNCONNECTED_45, SYNOPSYS_UNCONNECTED_46, 
        SYNOPSYS_UNCONNECTED_47, SYNOPSYS_UNCONNECTED_48, 
        SYNOPSYS_UNCONNECTED_49, SYNOPSYS_UNCONNECTED_50, 
        SYNOPSYS_UNCONNECTED_51, SYNOPSYS_UNCONNECTED_52, 
        SYNOPSYS_UNCONNECTED_53, SYNOPSYS_UNCONNECTED_54, 
        SYNOPSYS_UNCONNECTED_55, SYNOPSYS_UNCONNECTED_56, 
        SYNOPSYS_UNCONNECTED_57, SYNOPSYS_UNCONNECTED_58, 
        SYNOPSYS_UNCONNECTED_59, SYNOPSYS_UNCONNECTED_60, 
        SYNOPSYS_UNCONNECTED_61, SYNOPSYS_UNCONNECTED_62, 
        SYNOPSYS_UNCONNECTED_63, SYNOPSYS_UNCONNECTED_64, 
        SYNOPSYS_UNCONNECTED_65, SYNOPSYS_UNCONNECTED_66, 
        SYNOPSYS_UNCONNECTED_67, SYNOPSYS_UNCONNECTED_68, 
        SYNOPSYS_UNCONNECTED_69, SYNOPSYS_UNCONNECTED_70, 
        SYNOPSYS_UNCONNECTED_71, SYNOPSYS_UNCONNECTED_72, 
        SYNOPSYS_UNCONNECTED_73, SYNOPSYS_UNCONNECTED_74, 
        SYNOPSYS_UNCONNECTED_75, SYNOPSYS_UNCONNECTED_76, 
        SYNOPSYS_UNCONNECTED_77, SYNOPSYS_UNCONNECTED_78, 
        SYNOPSYS_UNCONNECTED_79, SYNOPSYS_UNCONNECTED_80, 
        SYNOPSYS_UNCONNECTED_81, SYNOPSYS_UNCONNECTED_82, 
        SYNOPSYS_UNCONNECTED_83, SYNOPSYS_UNCONNECTED_84, 
        SYNOPSYS_UNCONNECTED_85, SYNOPSYS_UNCONNECTED_86, 
        SYNOPSYS_UNCONNECTED_87, SYNOPSYS_UNCONNECTED_88, 
        SYNOPSYS_UNCONNECTED_89, SYNOPSYS_UNCONNECTED_90, 
        SYNOPSYS_UNCONNECTED_91, SYNOPSYS_UNCONNECTED_92, 
        SYNOPSYS_UNCONNECTED_93, SYNOPSYS_UNCONNECTED_94, 
        SYNOPSYS_UNCONNECTED_95, SYNOPSYS_UNCONNECTED_96, 
        SYNOPSYS_UNCONNECTED_97, SYNOPSYS_UNCONNECTED_98, 
        SYNOPSYS_UNCONNECTED_99, SYNOPSYS_UNCONNECTED_100, 
        SYNOPSYS_UNCONNECTED_101, SYNOPSYS_UNCONNECTED_102, 
        SYNOPSYS_UNCONNECTED_103, SYNOPSYS_UNCONNECTED_104, 
        SYNOPSYS_UNCONNECTED_105, SYNOPSYS_UNCONNECTED_106, 
        SYNOPSYS_UNCONNECTED_107, SYNOPSYS_UNCONNECTED_108, 
        SYNOPSYS_UNCONNECTED_109, SYNOPSYS_UNCONNECTED_110, 
        SYNOPSYS_UNCONNECTED_111, SYNOPSYS_UNCONNECTED_112, 
        SYNOPSYS_UNCONNECTED_113, SYNOPSYS_UNCONNECTED_114, 
        SYNOPSYS_UNCONNECTED_115, SYNOPSYS_UNCONNECTED_116, 
        SYNOPSYS_UNCONNECTED_117, SYNOPSYS_UNCONNECTED_118, 
        SYNOPSYS_UNCONNECTED_119, SYNOPSYS_UNCONNECTED_120, 
        SYNOPSYS_UNCONNECTED_121, SYNOPSYS_UNCONNECTED_122, 
        SYNOPSYS_UNCONNECTED_123, SYNOPSYS_UNCONNECTED_124, 
        SYNOPSYS_UNCONNECTED_125, SYNOPSYS_UNCONNECTED_126, 
        SYNOPSYS_UNCONNECTED_127, SYNOPSYS_UNCONNECTED_128, 
        SYNOPSYS_UNCONNECTED_129, SYNOPSYS_UNCONNECTED_130, 
        SYNOPSYS_UNCONNECTED_131, SYNOPSYS_UNCONNECTED_132, 
        SYNOPSYS_UNCONNECTED_133, SYNOPSYS_UNCONNECTED_134, 
        SYNOPSYS_UNCONNECTED_135, SYNOPSYS_UNCONNECTED_136, 
        SYNOPSYS_UNCONNECTED_137, SYNOPSYS_UNCONNECTED_138, 
        SYNOPSYS_UNCONNECTED_139, SYNOPSYS_UNCONNECTED_140, 
        SYNOPSYS_UNCONNECTED_141, SYNOPSYS_UNCONNECTED_142, 
        SYNOPSYS_UNCONNECTED_143, SYNOPSYS_UNCONNECTED_144, 
        SYNOPSYS_UNCONNECTED_145, SYNOPSYS_UNCONNECTED_146, 
        SYNOPSYS_UNCONNECTED_147, SYNOPSYS_UNCONNECTED_148, 
        SYNOPSYS_UNCONNECTED_149, SYNOPSYS_UNCONNECTED_150, 
        SYNOPSYS_UNCONNECTED_151, SYNOPSYS_UNCONNECTED_152, 
        SYNOPSYS_UNCONNECTED_153, SYNOPSYS_UNCONNECTED_154, 
        SYNOPSYS_UNCONNECTED_155, SYNOPSYS_UNCONNECTED_156, 
        SYNOPSYS_UNCONNECTED_157, SYNOPSYS_UNCONNECTED_158, 
        SYNOPSYS_UNCONNECTED_159, SYNOPSYS_UNCONNECTED_160, 
        SYNOPSYS_UNCONNECTED_161, SYNOPSYS_UNCONNECTED_162, 
        SYNOPSYS_UNCONNECTED_163, SYNOPSYS_UNCONNECTED_164, 
        SYNOPSYS_UNCONNECTED_165, SYNOPSYS_UNCONNECTED_166, 
        SYNOPSYS_UNCONNECTED_167, SYNOPSYS_UNCONNECTED_168, 
        SYNOPSYS_UNCONNECTED_169, SYNOPSYS_UNCONNECTED_170, 
        SYNOPSYS_UNCONNECTED_171, SYNOPSYS_UNCONNECTED_172, 
        SYNOPSYS_UNCONNECTED_173, SYNOPSYS_UNCONNECTED_174, 
        SYNOPSYS_UNCONNECTED_175, SYNOPSYS_UNCONNECTED_176, 
        SYNOPSYS_UNCONNECTED_177, SYNOPSYS_UNCONNECTED_178, 
        SYNOPSYS_UNCONNECTED_179, SYNOPSYS_UNCONNECTED_180, 
        SYNOPSYS_UNCONNECTED_181, SYNOPSYS_UNCONNECTED_182, 
        SYNOPSYS_UNCONNECTED_183, SYNOPSYS_UNCONNECTED_184, 
        SYNOPSYS_UNCONNECTED_185, SYNOPSYS_UNCONNECTED_186, 
        SYNOPSYS_UNCONNECTED_187, SYNOPSYS_UNCONNECTED_188, 
        SYNOPSYS_UNCONNECTED_189, SYNOPSYS_UNCONNECTED_190, 
        SYNOPSYS_UNCONNECTED_191, SYNOPSYS_UNCONNECTED_192, 
        SYNOPSYS_UNCONNECTED_193, SYNOPSYS_UNCONNECTED_194, 
        SYNOPSYS_UNCONNECTED_195, SYNOPSYS_UNCONNECTED_196, 
        SYNOPSYS_UNCONNECTED_197, SYNOPSYS_UNCONNECTED_198, 
        SYNOPSYS_UNCONNECTED_199, SYNOPSYS_UNCONNECTED_200, 
        SYNOPSYS_UNCONNECTED_201, SYNOPSYS_UNCONNECTED_202, 
        SYNOPSYS_UNCONNECTED_203, SYNOPSYS_UNCONNECTED_204, 
        SYNOPSYS_UNCONNECTED_205, SYNOPSYS_UNCONNECTED_206, 
        SYNOPSYS_UNCONNECTED_207, SYNOPSYS_UNCONNECTED_208, 
        SYNOPSYS_UNCONNECTED_209, SYNOPSYS_UNCONNECTED_210, 
        SYNOPSYS_UNCONNECTED_211, SYNOPSYS_UNCONNECTED_212, 
        SYNOPSYS_UNCONNECTED_213, SYNOPSYS_UNCONNECTED_214, 
        SYNOPSYS_UNCONNECTED_215, SYNOPSYS_UNCONNECTED_216, 
        SYNOPSYS_UNCONNECTED_217, SYNOPSYS_UNCONNECTED_218, 
        SYNOPSYS_UNCONNECTED_219, SYNOPSYS_UNCONNECTED_220, 
        SYNOPSYS_UNCONNECTED_221, SYNOPSYS_UNCONNECTED_222, 
        SYNOPSYS_UNCONNECTED_223, SYNOPSYS_UNCONNECTED_224, 
        SYNOPSYS_UNCONNECTED_225, SYNOPSYS_UNCONNECTED_226, 
        SYNOPSYS_UNCONNECTED_227, SYNOPSYS_UNCONNECTED_228, 
        SYNOPSYS_UNCONNECTED_229, SYNOPSYS_UNCONNECTED_230, 
        SYNOPSYS_UNCONNECTED_231, SYNOPSYS_UNCONNECTED_232, 
        SYNOPSYS_UNCONNECTED_233, SYNOPSYS_UNCONNECTED_234, 
        SYNOPSYS_UNCONNECTED_235, SYNOPSYS_UNCONNECTED_236, 
        SYNOPSYS_UNCONNECTED_237, SYNOPSYS_UNCONNECTED_238, 
        SYNOPSYS_UNCONNECTED_239, SYNOPSYS_UNCONNECTED_240, 
        SYNOPSYS_UNCONNECTED_241, SYNOPSYS_UNCONNECTED_242, 
        SYNOPSYS_UNCONNECTED_243, SYNOPSYS_UNCONNECTED_244, 
        SYNOPSYS_UNCONNECTED_245, SYNOPSYS_UNCONNECTED_246, 
        SYNOPSYS_UNCONNECTED_247, SYNOPSYS_UNCONNECTED_248, 
        SYNOPSYS_UNCONNECTED_249, SYNOPSYS_UNCONNECTED_250, 
        SYNOPSYS_UNCONNECTED_251, SYNOPSYS_UNCONNECTED_252, 
        SYNOPSYS_UNCONNECTED_253, SYNOPSYS_UNCONNECTED_254, 
        SYNOPSYS_UNCONNECTED_255, SYNOPSYS_UNCONNECTED_256, 
        SYNOPSYS_UNCONNECTED_257, SYNOPSYS_UNCONNECTED_258, 
        SYNOPSYS_UNCONNECTED_259, SYNOPSYS_UNCONNECTED_260, 
        SYNOPSYS_UNCONNECTED_261, SYNOPSYS_UNCONNECTED_262, 
        SYNOPSYS_UNCONNECTED_263, SYNOPSYS_UNCONNECTED_264, 
        SYNOPSYS_UNCONNECTED_265, SYNOPSYS_UNCONNECTED_266, 
        SYNOPSYS_UNCONNECTED_267, SYNOPSYS_UNCONNECTED_268, 
        SYNOPSYS_UNCONNECTED_269, SYNOPSYS_UNCONNECTED_270, 
        SYNOPSYS_UNCONNECTED_271, SYNOPSYS_UNCONNECTED_272, 
        SYNOPSYS_UNCONNECTED_273, SYNOPSYS_UNCONNECTED_274, 
        SYNOPSYS_UNCONNECTED_275, SYNOPSYS_UNCONNECTED_276, 
        SYNOPSYS_UNCONNECTED_277, SYNOPSYS_UNCONNECTED_278, 
        SYNOPSYS_UNCONNECTED_279, SYNOPSYS_UNCONNECTED_280, 
        SYNOPSYS_UNCONNECTED_281, SYNOPSYS_UNCONNECTED_282, 
        SYNOPSYS_UNCONNECTED_283, SYNOPSYS_UNCONNECTED_284, 
        SYNOPSYS_UNCONNECTED_285, SYNOPSYS_UNCONNECTED_286, 
        SYNOPSYS_UNCONNECTED_287, SYNOPSYS_UNCONNECTED_288, 
        SYNOPSYS_UNCONNECTED_289, SYNOPSYS_UNCONNECTED_290, 
        SYNOPSYS_UNCONNECTED_291, SYNOPSYS_UNCONNECTED_292, 
        SYNOPSYS_UNCONNECTED_293, SYNOPSYS_UNCONNECTED_294, 
        SYNOPSYS_UNCONNECTED_295, SYNOPSYS_UNCONNECTED_296, 
        SYNOPSYS_UNCONNECTED_297, SYNOPSYS_UNCONNECTED_298, 
        SYNOPSYS_UNCONNECTED_299, SYNOPSYS_UNCONNECTED_300, 
        SYNOPSYS_UNCONNECTED_301, SYNOPSYS_UNCONNECTED_302, 
        SYNOPSYS_UNCONNECTED_303, SYNOPSYS_UNCONNECTED_304, 
        SYNOPSYS_UNCONNECTED_305, SYNOPSYS_UNCONNECTED_306, 
        SYNOPSYS_UNCONNECTED_307, SYNOPSYS_UNCONNECTED_308, 
        SYNOPSYS_UNCONNECTED_309, SYNOPSYS_UNCONNECTED_310, 
        SYNOPSYS_UNCONNECTED_311, SYNOPSYS_UNCONNECTED_312, 
        SYNOPSYS_UNCONNECTED_313, SYNOPSYS_UNCONNECTED_314, 
        SYNOPSYS_UNCONNECTED_315, SYNOPSYS_UNCONNECTED_316, 
        SYNOPSYS_UNCONNECTED_317, SYNOPSYS_UNCONNECTED_318, 
        SYNOPSYS_UNCONNECTED_319, SYNOPSYS_UNCONNECTED_320, 
        SYNOPSYS_UNCONNECTED_321, SYNOPSYS_UNCONNECTED_322, 
        SYNOPSYS_UNCONNECTED_323, SYNOPSYS_UNCONNECTED_324, 
        SYNOPSYS_UNCONNECTED_325, SYNOPSYS_UNCONNECTED_326, 
        SYNOPSYS_UNCONNECTED_327, SYNOPSYS_UNCONNECTED_328, 
        SYNOPSYS_UNCONNECTED_329, SYNOPSYS_UNCONNECTED_330, 
        SYNOPSYS_UNCONNECTED_331, SYNOPSYS_UNCONNECTED_332, 
        SYNOPSYS_UNCONNECTED_333, SYNOPSYS_UNCONNECTED_334, 
        SYNOPSYS_UNCONNECTED_335, SYNOPSYS_UNCONNECTED_336, 
        SYNOPSYS_UNCONNECTED_337, SYNOPSYS_UNCONNECTED_338, 
        SYNOPSYS_UNCONNECTED_339, SYNOPSYS_UNCONNECTED_340, 
        SYNOPSYS_UNCONNECTED_341, SYNOPSYS_UNCONNECTED_342, 
        SYNOPSYS_UNCONNECTED_343, SYNOPSYS_UNCONNECTED_344, 
        SYNOPSYS_UNCONNECTED_345, SYNOPSYS_UNCONNECTED_346, 
        SYNOPSYS_UNCONNECTED_347, SYNOPSYS_UNCONNECTED_348, 
        SYNOPSYS_UNCONNECTED_349, SYNOPSYS_UNCONNECTED_350, 
        SYNOPSYS_UNCONNECTED_351, SYNOPSYS_UNCONNECTED_352, 
        SYNOPSYS_UNCONNECTED_353, SYNOPSYS_UNCONNECTED_354, 
        SYNOPSYS_UNCONNECTED_355, SYNOPSYS_UNCONNECTED_356, 
        SYNOPSYS_UNCONNECTED_357, SYNOPSYS_UNCONNECTED_358, 
        SYNOPSYS_UNCONNECTED_359, SYNOPSYS_UNCONNECTED_360, 
        SYNOPSYS_UNCONNECTED_361, SYNOPSYS_UNCONNECTED_362, 
        SYNOPSYS_UNCONNECTED_363, SYNOPSYS_UNCONNECTED_364, 
        SYNOPSYS_UNCONNECTED_365, SYNOPSYS_UNCONNECTED_366, 
        SYNOPSYS_UNCONNECTED_367, SYNOPSYS_UNCONNECTED_368, 
        SYNOPSYS_UNCONNECTED_369, SYNOPSYS_UNCONNECTED_370, 
        SYNOPSYS_UNCONNECTED_371, SYNOPSYS_UNCONNECTED_372, 
        SYNOPSYS_UNCONNECTED_373, SYNOPSYS_UNCONNECTED_374, 
        SYNOPSYS_UNCONNECTED_375, SYNOPSYS_UNCONNECTED_376, 
        SYNOPSYS_UNCONNECTED_377, SYNOPSYS_UNCONNECTED_378, 
        SYNOPSYS_UNCONNECTED_379, SYNOPSYS_UNCONNECTED_380, 
        SYNOPSYS_UNCONNECTED_381, SYNOPSYS_UNCONNECTED_382, 
        SYNOPSYS_UNCONNECTED_383, SYNOPSYS_UNCONNECTED_384, 
        SYNOPSYS_UNCONNECTED_385, SYNOPSYS_UNCONNECTED_386, 
        SYNOPSYS_UNCONNECTED_387, SYNOPSYS_UNCONNECTED_388, 
        SYNOPSYS_UNCONNECTED_389, SYNOPSYS_UNCONNECTED_390, 
        SYNOPSYS_UNCONNECTED_391, SYNOPSYS_UNCONNECTED_392, 
        SYNOPSYS_UNCONNECTED_393, SYNOPSYS_UNCONNECTED_394, 
        SYNOPSYS_UNCONNECTED_395, SYNOPSYS_UNCONNECTED_396, 
        SYNOPSYS_UNCONNECTED_397, SYNOPSYS_UNCONNECTED_398, 
        SYNOPSYS_UNCONNECTED_399, SYNOPSYS_UNCONNECTED_400, 
        SYNOPSYS_UNCONNECTED_401, SYNOPSYS_UNCONNECTED_402, 
        SYNOPSYS_UNCONNECTED_403, SYNOPSYS_UNCONNECTED_404, 
        SYNOPSYS_UNCONNECTED_405, SYNOPSYS_UNCONNECTED_406, 
        SYNOPSYS_UNCONNECTED_407, SYNOPSYS_UNCONNECTED_408, 
        SYNOPSYS_UNCONNECTED_409, SYNOPSYS_UNCONNECTED_410, 
        SYNOPSYS_UNCONNECTED_411, SYNOPSYS_UNCONNECTED_412, 
        SYNOPSYS_UNCONNECTED_413, SYNOPSYS_UNCONNECTED_414, 
        SYNOPSYS_UNCONNECTED_415, SYNOPSYS_UNCONNECTED_416, 
        SYNOPSYS_UNCONNECTED_417, SYNOPSYS_UNCONNECTED_418, 
        SYNOPSYS_UNCONNECTED_419, SYNOPSYS_UNCONNECTED_420, 
        SYNOPSYS_UNCONNECTED_421, SYNOPSYS_UNCONNECTED_422, 
        SYNOPSYS_UNCONNECTED_423, SYNOPSYS_UNCONNECTED_424, 
        SYNOPSYS_UNCONNECTED_425, SYNOPSYS_UNCONNECTED_426, 
        SYNOPSYS_UNCONNECTED_427, SYNOPSYS_UNCONNECTED_428, 
        SYNOPSYS_UNCONNECTED_429, SYNOPSYS_UNCONNECTED_430, 
        SYNOPSYS_UNCONNECTED_431, SYNOPSYS_UNCONNECTED_432, 
        SYNOPSYS_UNCONNECTED_433, SYNOPSYS_UNCONNECTED_434, 
        SYNOPSYS_UNCONNECTED_435, SYNOPSYS_UNCONNECTED_436, 
        SYNOPSYS_UNCONNECTED_437, SYNOPSYS_UNCONNECTED_438, 
        SYNOPSYS_UNCONNECTED_439, SYNOPSYS_UNCONNECTED_440, 
        SYNOPSYS_UNCONNECTED_441, SYNOPSYS_UNCONNECTED_442, 
        SYNOPSYS_UNCONNECTED_443, SYNOPSYS_UNCONNECTED_444, 
        SYNOPSYS_UNCONNECTED_445, SYNOPSYS_UNCONNECTED_446, 
        SYNOPSYS_UNCONNECTED_447, SYNOPSYS_UNCONNECTED_448, 
        SYNOPSYS_UNCONNECTED_449, SYNOPSYS_UNCONNECTED_450, 
        SYNOPSYS_UNCONNECTED_451, SYNOPSYS_UNCONNECTED_452, 
        SYNOPSYS_UNCONNECTED_453, SYNOPSYS_UNCONNECTED_454, 
        SYNOPSYS_UNCONNECTED_455, SYNOPSYS_UNCONNECTED_456, 
        SYNOPSYS_UNCONNECTED_457, SYNOPSYS_UNCONNECTED_458, 
        SYNOPSYS_UNCONNECTED_459, SYNOPSYS_UNCONNECTED_460, 
        SYNOPSYS_UNCONNECTED_461, SYNOPSYS_UNCONNECTED_462, 
        SYNOPSYS_UNCONNECTED_463, SYNOPSYS_UNCONNECTED_464, 
        SYNOPSYS_UNCONNECTED_465, SYNOPSYS_UNCONNECTED_466, 
        SYNOPSYS_UNCONNECTED_467, SYNOPSYS_UNCONNECTED_468, 
        SYNOPSYS_UNCONNECTED_469, SYNOPSYS_UNCONNECTED_470, 
        SYNOPSYS_UNCONNECTED_471, SYNOPSYS_UNCONNECTED_472, 
        SYNOPSYS_UNCONNECTED_473, SYNOPSYS_UNCONNECTED_474, 
        SYNOPSYS_UNCONNECTED_475, SYNOPSYS_UNCONNECTED_476, 
        SYNOPSYS_UNCONNECTED_477, SYNOPSYS_UNCONNECTED_478, 
        SYNOPSYS_UNCONNECTED_479, SYNOPSYS_UNCONNECTED_480, 
        SYNOPSYS_UNCONNECTED_481, SYNOPSYS_UNCONNECTED_482, 
        SYNOPSYS_UNCONNECTED_483, SYNOPSYS_UNCONNECTED_484, 
        SYNOPSYS_UNCONNECTED_485, SYNOPSYS_UNCONNECTED_486, 
        SYNOPSYS_UNCONNECTED_487, SYNOPSYS_UNCONNECTED_488, 
        SYNOPSYS_UNCONNECTED_489, SYNOPSYS_UNCONNECTED_490, 
        SYNOPSYS_UNCONNECTED_491, SYNOPSYS_UNCONNECTED_492, 
        SYNOPSYS_UNCONNECTED_493, SYNOPSYS_UNCONNECTED_494, 
        SYNOPSYS_UNCONNECTED_495, SYNOPSYS_UNCONNECTED_496, 
        SYNOPSYS_UNCONNECTED_497, SYNOPSYS_UNCONNECTED_498, 
        SYNOPSYS_UNCONNECTED_499, SYNOPSYS_UNCONNECTED_500, 
        SYNOPSYS_UNCONNECTED_501, SYNOPSYS_UNCONNECTED_502, 
        SYNOPSYS_UNCONNECTED_503, SYNOPSYS_UNCONNECTED_504, 
        SYNOPSYS_UNCONNECTED_505, SYNOPSYS_UNCONNECTED_506, 
        SYNOPSYS_UNCONNECTED_507, SYNOPSYS_UNCONNECTED_508, 
        SYNOPSYS_UNCONNECTED_509, SYNOPSYS_UNCONNECTED_510, 
        SYNOPSYS_UNCONNECTED_511, SYNOPSYS_UNCONNECTED_512, 
        SYNOPSYS_UNCONNECTED_513, SYNOPSYS_UNCONNECTED_514, 
        SYNOPSYS_UNCONNECTED_515, SYNOPSYS_UNCONNECTED_516, 
        SYNOPSYS_UNCONNECTED_517, SYNOPSYS_UNCONNECTED_518, 
        SYNOPSYS_UNCONNECTED_519, SYNOPSYS_UNCONNECTED_520, 
        SYNOPSYS_UNCONNECTED_521, SYNOPSYS_UNCONNECTED_522, 
        SYNOPSYS_UNCONNECTED_523, SYNOPSYS_UNCONNECTED_524, 
        SYNOPSYS_UNCONNECTED_525, SYNOPSYS_UNCONNECTED_526, 
        SYNOPSYS_UNCONNECTED_527, SYNOPSYS_UNCONNECTED_528, 
        SYNOPSYS_UNCONNECTED_529, SYNOPSYS_UNCONNECTED_530, 
        SYNOPSYS_UNCONNECTED_531, SYNOPSYS_UNCONNECTED_532, 
        SYNOPSYS_UNCONNECTED_533, SYNOPSYS_UNCONNECTED_534, 
        SYNOPSYS_UNCONNECTED_535, SYNOPSYS_UNCONNECTED_536, 
        SYNOPSYS_UNCONNECTED_537, SYNOPSYS_UNCONNECTED_538, 
        SYNOPSYS_UNCONNECTED_539, SYNOPSYS_UNCONNECTED_540, 
        SYNOPSYS_UNCONNECTED_541, SYNOPSYS_UNCONNECTED_542, 
        SYNOPSYS_UNCONNECTED_543, SYNOPSYS_UNCONNECTED_544, 
        SYNOPSYS_UNCONNECTED_545, SYNOPSYS_UNCONNECTED_546, 
        SYNOPSYS_UNCONNECTED_547, SYNOPSYS_UNCONNECTED_548, 
        SYNOPSYS_UNCONNECTED_549, SYNOPSYS_UNCONNECTED_550, 
        SYNOPSYS_UNCONNECTED_551, SYNOPSYS_UNCONNECTED_552, 
        SYNOPSYS_UNCONNECTED_553, SYNOPSYS_UNCONNECTED_554, 
        SYNOPSYS_UNCONNECTED_555, SYNOPSYS_UNCONNECTED_556, 
        SYNOPSYS_UNCONNECTED_557, SYNOPSYS_UNCONNECTED_558, 
        SYNOPSYS_UNCONNECTED_559, SYNOPSYS_UNCONNECTED_560, 
        SYNOPSYS_UNCONNECTED_561, SYNOPSYS_UNCONNECTED_562, 
        SYNOPSYS_UNCONNECTED_563, SYNOPSYS_UNCONNECTED_564, 
        SYNOPSYS_UNCONNECTED_565, SYNOPSYS_UNCONNECTED_566, 
        SYNOPSYS_UNCONNECTED_567, SYNOPSYS_UNCONNECTED_568, 
        SYNOPSYS_UNCONNECTED_569, SYNOPSYS_UNCONNECTED_570, 
        SYNOPSYS_UNCONNECTED_571, SYNOPSYS_UNCONNECTED_572, 
        SYNOPSYS_UNCONNECTED_573, SYNOPSYS_UNCONNECTED_574, 
        SYNOPSYS_UNCONNECTED_575, SYNOPSYS_UNCONNECTED_576, 
        SYNOPSYS_UNCONNECTED_577, SYNOPSYS_UNCONNECTED_578, 
        SYNOPSYS_UNCONNECTED_579, SYNOPSYS_UNCONNECTED_580, 
        SYNOPSYS_UNCONNECTED_581, SYNOPSYS_UNCONNECTED_582, 
        SYNOPSYS_UNCONNECTED_583, SYNOPSYS_UNCONNECTED_584, 
        SYNOPSYS_UNCONNECTED_585, SYNOPSYS_UNCONNECTED_586, 
        SYNOPSYS_UNCONNECTED_587, SYNOPSYS_UNCONNECTED_588, 
        SYNOPSYS_UNCONNECTED_589, SYNOPSYS_UNCONNECTED_590, 
        SYNOPSYS_UNCONNECTED_591, SYNOPSYS_UNCONNECTED_592, 
        SYNOPSYS_UNCONNECTED_593, SYNOPSYS_UNCONNECTED_594, 
        SYNOPSYS_UNCONNECTED_595, SYNOPSYS_UNCONNECTED_596, 
        SYNOPSYS_UNCONNECTED_597, SYNOPSYS_UNCONNECTED_598, 
        SYNOPSYS_UNCONNECTED_599, SYNOPSYS_UNCONNECTED_600, 
        SYNOPSYS_UNCONNECTED_601, SYNOPSYS_UNCONNECTED_602, 
        SYNOPSYS_UNCONNECTED_603, SYNOPSYS_UNCONNECTED_604, 
        SYNOPSYS_UNCONNECTED_605, SYNOPSYS_UNCONNECTED_606, 
        SYNOPSYS_UNCONNECTED_607, SYNOPSYS_UNCONNECTED_608, 
        SYNOPSYS_UNCONNECTED_609, SYNOPSYS_UNCONNECTED_610, 
        SYNOPSYS_UNCONNECTED_611, SYNOPSYS_UNCONNECTED_612, 
        SYNOPSYS_UNCONNECTED_613, SYNOPSYS_UNCONNECTED_614, 
        SYNOPSYS_UNCONNECTED_615, SYNOPSYS_UNCONNECTED_616, 
        SYNOPSYS_UNCONNECTED_617, SYNOPSYS_UNCONNECTED_618, 
        SYNOPSYS_UNCONNECTED_619, SYNOPSYS_UNCONNECTED_620, 
        SYNOPSYS_UNCONNECTED_621, SYNOPSYS_UNCONNECTED_622, 
        SYNOPSYS_UNCONNECTED_623, SYNOPSYS_UNCONNECTED_624, 
        SYNOPSYS_UNCONNECTED_625, SYNOPSYS_UNCONNECTED_626, 
        SYNOPSYS_UNCONNECTED_627, SYNOPSYS_UNCONNECTED_628, 
        SYNOPSYS_UNCONNECTED_629, SYNOPSYS_UNCONNECTED_630, 
        SYNOPSYS_UNCONNECTED_631, SYNOPSYS_UNCONNECTED_632, 
        SYNOPSYS_UNCONNECTED_633, SYNOPSYS_UNCONNECTED_634, 
        SYNOPSYS_UNCONNECTED_635, SYNOPSYS_UNCONNECTED_636, 
        SYNOPSYS_UNCONNECTED_637, SYNOPSYS_UNCONNECTED_638, 
        SYNOPSYS_UNCONNECTED_639, SYNOPSYS_UNCONNECTED_640, 
        SYNOPSYS_UNCONNECTED_641, SYNOPSYS_UNCONNECTED_642, 
        SYNOPSYS_UNCONNECTED_643, SYNOPSYS_UNCONNECTED_644, 
        SYNOPSYS_UNCONNECTED_645, SYNOPSYS_UNCONNECTED_646, 
        SYNOPSYS_UNCONNECTED_647, SYNOPSYS_UNCONNECTED_648, 
        SYNOPSYS_UNCONNECTED_649, SYNOPSYS_UNCONNECTED_650, 
        SYNOPSYS_UNCONNECTED_651, SYNOPSYS_UNCONNECTED_652, 
        SYNOPSYS_UNCONNECTED_653, SYNOPSYS_UNCONNECTED_654, 
        SYNOPSYS_UNCONNECTED_655, SYNOPSYS_UNCONNECTED_656, 
        SYNOPSYS_UNCONNECTED_657, SYNOPSYS_UNCONNECTED_658, 
        SYNOPSYS_UNCONNECTED_659, SYNOPSYS_UNCONNECTED_660, 
        SYNOPSYS_UNCONNECTED_661, SYNOPSYS_UNCONNECTED_662, 
        SYNOPSYS_UNCONNECTED_663, SYNOPSYS_UNCONNECTED_664, 
        SYNOPSYS_UNCONNECTED_665, SYNOPSYS_UNCONNECTED_666, 
        SYNOPSYS_UNCONNECTED_667, SYNOPSYS_UNCONNECTED_668, 
        SYNOPSYS_UNCONNECTED_669, SYNOPSYS_UNCONNECTED_670, 
        SYNOPSYS_UNCONNECTED_671, SYNOPSYS_UNCONNECTED_672, 
        SYNOPSYS_UNCONNECTED_673, SYNOPSYS_UNCONNECTED_674, 
        SYNOPSYS_UNCONNECTED_675, SYNOPSYS_UNCONNECTED_676, 
        SYNOPSYS_UNCONNECTED_677, SYNOPSYS_UNCONNECTED_678, 
        SYNOPSYS_UNCONNECTED_679, SYNOPSYS_UNCONNECTED_680, 
        SYNOPSYS_UNCONNECTED_681, SYNOPSYS_UNCONNECTED_682, 
        SYNOPSYS_UNCONNECTED_683, SYNOPSYS_UNCONNECTED_684, 
        SYNOPSYS_UNCONNECTED_685, SYNOPSYS_UNCONNECTED_686, 
        SYNOPSYS_UNCONNECTED_687, SYNOPSYS_UNCONNECTED_688, 
        SYNOPSYS_UNCONNECTED_689, SYNOPSYS_UNCONNECTED_690, 
        SYNOPSYS_UNCONNECTED_691, SYNOPSYS_UNCONNECTED_692, 
        SYNOPSYS_UNCONNECTED_693, SYNOPSYS_UNCONNECTED_694, 
        SYNOPSYS_UNCONNECTED_695, SYNOPSYS_UNCONNECTED_696, 
        SYNOPSYS_UNCONNECTED_697, SYNOPSYS_UNCONNECTED_698, 
        SYNOPSYS_UNCONNECTED_699, SYNOPSYS_UNCONNECTED_700, 
        SYNOPSYS_UNCONNECTED_701, SYNOPSYS_UNCONNECTED_702, 
        SYNOPSYS_UNCONNECTED_703, SYNOPSYS_UNCONNECTED_704, 
        SYNOPSYS_UNCONNECTED_705, SYNOPSYS_UNCONNECTED_706, 
        SYNOPSYS_UNCONNECTED_707, SYNOPSYS_UNCONNECTED_708, 
        SYNOPSYS_UNCONNECTED_709, SYNOPSYS_UNCONNECTED_710, 
        SYNOPSYS_UNCONNECTED_711, SYNOPSYS_UNCONNECTED_712, 
        SYNOPSYS_UNCONNECTED_713, SYNOPSYS_UNCONNECTED_714, 
        SYNOPSYS_UNCONNECTED_715, SYNOPSYS_UNCONNECTED_716, 
        SYNOPSYS_UNCONNECTED_717, SYNOPSYS_UNCONNECTED_718, 
        SYNOPSYS_UNCONNECTED_719, SYNOPSYS_UNCONNECTED_720, 
        SYNOPSYS_UNCONNECTED_721, SYNOPSYS_UNCONNECTED_722, 
        SYNOPSYS_UNCONNECTED_723, SYNOPSYS_UNCONNECTED_724, 
        SYNOPSYS_UNCONNECTED_725, SYNOPSYS_UNCONNECTED_726, 
        SYNOPSYS_UNCONNECTED_727, SYNOPSYS_UNCONNECTED_728, 
        SYNOPSYS_UNCONNECTED_729, SYNOPSYS_UNCONNECTED_730, 
        SYNOPSYS_UNCONNECTED_731, SYNOPSYS_UNCONNECTED_732, 
        SYNOPSYS_UNCONNECTED_733, SYNOPSYS_UNCONNECTED_734, 
        SYNOPSYS_UNCONNECTED_735, SYNOPSYS_UNCONNECTED_736, 
        SYNOPSYS_UNCONNECTED_737, SYNOPSYS_UNCONNECTED_738, 
        SYNOPSYS_UNCONNECTED_739, SYNOPSYS_UNCONNECTED_740, 
        SYNOPSYS_UNCONNECTED_741, SYNOPSYS_UNCONNECTED_742, 
        SYNOPSYS_UNCONNECTED_743, SYNOPSYS_UNCONNECTED_744, 
        SYNOPSYS_UNCONNECTED_745, SYNOPSYS_UNCONNECTED_746, 
        SYNOPSYS_UNCONNECTED_747, SYNOPSYS_UNCONNECTED_748, 
        SYNOPSYS_UNCONNECTED_749, SYNOPSYS_UNCONNECTED_750, 
        SYNOPSYS_UNCONNECTED_751, SYNOPSYS_UNCONNECTED_752, 
        SYNOPSYS_UNCONNECTED_753, SYNOPSYS_UNCONNECTED_754, 
        SYNOPSYS_UNCONNECTED_755, SYNOPSYS_UNCONNECTED_756, 
        SYNOPSYS_UNCONNECTED_757, SYNOPSYS_UNCONNECTED_758, 
        SYNOPSYS_UNCONNECTED_759, SYNOPSYS_UNCONNECTED_760, 
        SYNOPSYS_UNCONNECTED_761, SYNOPSYS_UNCONNECTED_762, 
        SYNOPSYS_UNCONNECTED_763, SYNOPSYS_UNCONNECTED_764, 
        SYNOPSYS_UNCONNECTED_765, SYNOPSYS_UNCONNECTED_766, 
        SYNOPSYS_UNCONNECTED_767, SYNOPSYS_UNCONNECTED_768, 
        SYNOPSYS_UNCONNECTED_769, SYNOPSYS_UNCONNECTED_770, 
        SYNOPSYS_UNCONNECTED_771, SYNOPSYS_UNCONNECTED_772, 
        SYNOPSYS_UNCONNECTED_773, SYNOPSYS_UNCONNECTED_774, 
        SYNOPSYS_UNCONNECTED_775, SYNOPSYS_UNCONNECTED_776, 
        SYNOPSYS_UNCONNECTED_777, SYNOPSYS_UNCONNECTED_778, 
        SYNOPSYS_UNCONNECTED_779, SYNOPSYS_UNCONNECTED_780, 
        SYNOPSYS_UNCONNECTED_781, SYNOPSYS_UNCONNECTED_782, 
        SYNOPSYS_UNCONNECTED_783, SYNOPSYS_UNCONNECTED_784, 
        SYNOPSYS_UNCONNECTED_785, SYNOPSYS_UNCONNECTED_786, 
        SYNOPSYS_UNCONNECTED_787, SYNOPSYS_UNCONNECTED_788, 
        SYNOPSYS_UNCONNECTED_789, SYNOPSYS_UNCONNECTED_790, 
        SYNOPSYS_UNCONNECTED_791, SYNOPSYS_UNCONNECTED_792, 
        SYNOPSYS_UNCONNECTED_793, SYNOPSYS_UNCONNECTED_794, 
        SYNOPSYS_UNCONNECTED_795, SYNOPSYS_UNCONNECTED_796, 
        SYNOPSYS_UNCONNECTED_797, SYNOPSYS_UNCONNECTED_798, 
        SYNOPSYS_UNCONNECTED_799, SYNOPSYS_UNCONNECTED_800, 
        SYNOPSYS_UNCONNECTED_801, SYNOPSYS_UNCONNECTED_802, 
        SYNOPSYS_UNCONNECTED_803, SYNOPSYS_UNCONNECTED_804, 
        SYNOPSYS_UNCONNECTED_805, SYNOPSYS_UNCONNECTED_806, 
        SYNOPSYS_UNCONNECTED_807, SYNOPSYS_UNCONNECTED_808, 
        SYNOPSYS_UNCONNECTED_809, SYNOPSYS_UNCONNECTED_810, 
        SYNOPSYS_UNCONNECTED_811, SYNOPSYS_UNCONNECTED_812, 
        SYNOPSYS_UNCONNECTED_813, SYNOPSYS_UNCONNECTED_814, 
        SYNOPSYS_UNCONNECTED_815, SYNOPSYS_UNCONNECTED_816, 
        SYNOPSYS_UNCONNECTED_817, SYNOPSYS_UNCONNECTED_818, 
        SYNOPSYS_UNCONNECTED_819, SYNOPSYS_UNCONNECTED_820, 
        SYNOPSYS_UNCONNECTED_821, SYNOPSYS_UNCONNECTED_822, 
        SYNOPSYS_UNCONNECTED_823, SYNOPSYS_UNCONNECTED_824, 
        SYNOPSYS_UNCONNECTED_825, SYNOPSYS_UNCONNECTED_826, 
        SYNOPSYS_UNCONNECTED_827, SYNOPSYS_UNCONNECTED_828, 
        SYNOPSYS_UNCONNECTED_829, SYNOPSYS_UNCONNECTED_830, 
        SYNOPSYS_UNCONNECTED_831, SYNOPSYS_UNCONNECTED_832, 
        SYNOPSYS_UNCONNECTED_833, SYNOPSYS_UNCONNECTED_834, 
        SYNOPSYS_UNCONNECTED_835, SYNOPSYS_UNCONNECTED_836, 
        SYNOPSYS_UNCONNECTED_837, SYNOPSYS_UNCONNECTED_838, 
        SYNOPSYS_UNCONNECTED_839, SYNOPSYS_UNCONNECTED_840, 
        SYNOPSYS_UNCONNECTED_841, SYNOPSYS_UNCONNECTED_842, 
        SYNOPSYS_UNCONNECTED_843, SYNOPSYS_UNCONNECTED_844, 
        SYNOPSYS_UNCONNECTED_845, SYNOPSYS_UNCONNECTED_846, 
        SYNOPSYS_UNCONNECTED_847, SYNOPSYS_UNCONNECTED_848, 
        SYNOPSYS_UNCONNECTED_849, SYNOPSYS_UNCONNECTED_850, 
        SYNOPSYS_UNCONNECTED_851, SYNOPSYS_UNCONNECTED_852, 
        SYNOPSYS_UNCONNECTED_853, SYNOPSYS_UNCONNECTED_854, 
        SYNOPSYS_UNCONNECTED_855, SYNOPSYS_UNCONNECTED_856, 
        SYNOPSYS_UNCONNECTED_857, SYNOPSYS_UNCONNECTED_858, 
        SYNOPSYS_UNCONNECTED_859, SYNOPSYS_UNCONNECTED_860, 
        SYNOPSYS_UNCONNECTED_861, SYNOPSYS_UNCONNECTED_862, 
        SYNOPSYS_UNCONNECTED_863, SYNOPSYS_UNCONNECTED_864, 
        SYNOPSYS_UNCONNECTED_865, SYNOPSYS_UNCONNECTED_866, 
        SYNOPSYS_UNCONNECTED_867, SYNOPSYS_UNCONNECTED_868, 
        SYNOPSYS_UNCONNECTED_869, SYNOPSYS_UNCONNECTED_870, 
        SYNOPSYS_UNCONNECTED_871, SYNOPSYS_UNCONNECTED_872, 
        SYNOPSYS_UNCONNECTED_873, SYNOPSYS_UNCONNECTED_874, 
        SYNOPSYS_UNCONNECTED_875, SYNOPSYS_UNCONNECTED_876, 
        SYNOPSYS_UNCONNECTED_877, SYNOPSYS_UNCONNECTED_878, 
        SYNOPSYS_UNCONNECTED_879, SYNOPSYS_UNCONNECTED_880, 
        SYNOPSYS_UNCONNECTED_881, SYNOPSYS_UNCONNECTED_882, 
        SYNOPSYS_UNCONNECTED_883, SYNOPSYS_UNCONNECTED_884, 
        SYNOPSYS_UNCONNECTED_885, SYNOPSYS_UNCONNECTED_886, 
        SYNOPSYS_UNCONNECTED_887, SYNOPSYS_UNCONNECTED_888, 
        SYNOPSYS_UNCONNECTED_889, SYNOPSYS_UNCONNECTED_890, 
        SYNOPSYS_UNCONNECTED_891, SYNOPSYS_UNCONNECTED_892, 
        SYNOPSYS_UNCONNECTED_893, SYNOPSYS_UNCONNECTED_894, 
        SYNOPSYS_UNCONNECTED_895, SYNOPSYS_UNCONNECTED_896, 
        SYNOPSYS_UNCONNECTED_897, SYNOPSYS_UNCONNECTED_898, 
        SYNOPSYS_UNCONNECTED_899, SYNOPSYS_UNCONNECTED_900, 
        SYNOPSYS_UNCONNECTED_901, SYNOPSYS_UNCONNECTED_902, 
        SYNOPSYS_UNCONNECTED_903, SYNOPSYS_UNCONNECTED_904, 
        SYNOPSYS_UNCONNECTED_905, SYNOPSYS_UNCONNECTED_906, 
        SYNOPSYS_UNCONNECTED_907, SYNOPSYS_UNCONNECTED_908, 
        SYNOPSYS_UNCONNECTED_909, SYNOPSYS_UNCONNECTED_910, 
        SYNOPSYS_UNCONNECTED_911, SYNOPSYS_UNCONNECTED_912, 
        SYNOPSYS_UNCONNECTED_913, SYNOPSYS_UNCONNECTED_914, 
        SYNOPSYS_UNCONNECTED_915, SYNOPSYS_UNCONNECTED_916, 
        SYNOPSYS_UNCONNECTED_917, SYNOPSYS_UNCONNECTED_918, 
        SYNOPSYS_UNCONNECTED_919, SYNOPSYS_UNCONNECTED_920, 
        SYNOPSYS_UNCONNECTED_921, SYNOPSYS_UNCONNECTED_922, 
        SYNOPSYS_UNCONNECTED_923, SYNOPSYS_UNCONNECTED_924, 
        SYNOPSYS_UNCONNECTED_925, SYNOPSYS_UNCONNECTED_926, 
        SYNOPSYS_UNCONNECTED_927, SYNOPSYS_UNCONNECTED_928, 
        SYNOPSYS_UNCONNECTED_929, SYNOPSYS_UNCONNECTED_930, 
        SYNOPSYS_UNCONNECTED_931, SYNOPSYS_UNCONNECTED_932, 
        SYNOPSYS_UNCONNECTED_933, SYNOPSYS_UNCONNECTED_934, 
        SYNOPSYS_UNCONNECTED_935, SYNOPSYS_UNCONNECTED_936, 
        SYNOPSYS_UNCONNECTED_937, SYNOPSYS_UNCONNECTED_938, 
        SYNOPSYS_UNCONNECTED_939, SYNOPSYS_UNCONNECTED_940, 
        SYNOPSYS_UNCONNECTED_941, SYNOPSYS_UNCONNECTED_942, 
        SYNOPSYS_UNCONNECTED_943, SYNOPSYS_UNCONNECTED_944, 
        SYNOPSYS_UNCONNECTED_945, SYNOPSYS_UNCONNECTED_946, 
        SYNOPSYS_UNCONNECTED_947, SYNOPSYS_UNCONNECTED_948, 
        SYNOPSYS_UNCONNECTED_949, SYNOPSYS_UNCONNECTED_950, 
        SYNOPSYS_UNCONNECTED_951, SYNOPSYS_UNCONNECTED_952, 
        SYNOPSYS_UNCONNECTED_953, SYNOPSYS_UNCONNECTED_954, 
        SYNOPSYS_UNCONNECTED_955, SYNOPSYS_UNCONNECTED_956, 
        SYNOPSYS_UNCONNECTED_957, SYNOPSYS_UNCONNECTED_958, 
        SYNOPSYS_UNCONNECTED_959, SYNOPSYS_UNCONNECTED_960, 
        SYNOPSYS_UNCONNECTED_961, SYNOPSYS_UNCONNECTED_962, 
        SYNOPSYS_UNCONNECTED_963, SYNOPSYS_UNCONNECTED_964, 
        SYNOPSYS_UNCONNECTED_965, SYNOPSYS_UNCONNECTED_966, 
        SYNOPSYS_UNCONNECTED_967, SYNOPSYS_UNCONNECTED_968, 
        SYNOPSYS_UNCONNECTED_969, SYNOPSYS_UNCONNECTED_970, 
        SYNOPSYS_UNCONNECTED_971, SYNOPSYS_UNCONNECTED_972, 
        SYNOPSYS_UNCONNECTED_973, SYNOPSYS_UNCONNECTED_974, 
        SYNOPSYS_UNCONNECTED_975, SYNOPSYS_UNCONNECTED_976, 
        SYNOPSYS_UNCONNECTED_977, SYNOPSYS_UNCONNECTED_978, 
        SYNOPSYS_UNCONNECTED_979, SYNOPSYS_UNCONNECTED_980, 
        SYNOPSYS_UNCONNECTED_981, SYNOPSYS_UNCONNECTED_982, 
        SYNOPSYS_UNCONNECTED_983, SYNOPSYS_UNCONNECTED_984, 
        SYNOPSYS_UNCONNECTED_985, SYNOPSYS_UNCONNECTED_986, 
        SYNOPSYS_UNCONNECTED_987, SYNOPSYS_UNCONNECTED_988, 
        SYNOPSYS_UNCONNECTED_989, SYNOPSYS_UNCONNECTED_990, 
        SYNOPSYS_UNCONNECTED_991, SYNOPSYS_UNCONNECTED_992, 
        SYNOPSYS_UNCONNECTED_993, SYNOPSYS_UNCONNECTED_994, 
        SYNOPSYS_UNCONNECTED_995, SYNOPSYS_UNCONNECTED_996, 
        SYNOPSYS_UNCONNECTED_997, SYNOPSYS_UNCONNECTED_998, 
        SYNOPSYS_UNCONNECTED_999, SYNOPSYS_UNCONNECTED_1000, 
        SYNOPSYS_UNCONNECTED_1001, SYNOPSYS_UNCONNECTED_1002, 
        SYNOPSYS_UNCONNECTED_1003, SYNOPSYS_UNCONNECTED_1004, 
        SYNOPSYS_UNCONNECTED_1005, SYNOPSYS_UNCONNECTED_1006, 
        SYNOPSYS_UNCONNECTED_1007, SYNOPSYS_UNCONNECTED_1008, 
        SYNOPSYS_UNCONNECTED_1009, SYNOPSYS_UNCONNECTED_1010, 
        SYNOPSYS_UNCONNECTED_1011, SYNOPSYS_UNCONNECTED_1012, 
        SYNOPSYS_UNCONNECTED_1013, SYNOPSYS_UNCONNECTED_1014, 
        SYNOPSYS_UNCONNECTED_1015, SYNOPSYS_UNCONNECTED_1016, regx_rdat}) );
  DFFQX1 d_regx_addr_reg_2_ ( .D(regx_addr[2]), .C(clk), .Q(d_regx_addr[2]) );
  DFFQX1 d_we16_reg ( .D(N8), .C(clk), .Q(d_we16) );
  DFFQX1 d_lt_drp_reg ( .D(lt_drp), .C(clk), .Q(reg14[0]) );
  DFFQX1 d_di_tst_reg ( .D(di_tst), .C(clk), .Q(reg14[3]) );
  DFFQX1 d_lt_gpi_reg_1_ ( .D(lt_gpi[1]), .C(net8975), .Q(d_lt_gpi[1]) );
  DFFQX1 d_lt_gpi_reg_0_ ( .D(lt_gpi[0]), .C(net8975), .Q(d_lt_gpi[0]) );
  DFFQX1 d_lt_aswk_reg_5_ ( .D(lt_aswk[5]), .C(clk), .Q(d_lt_aswk[5]) );
  DFFQX1 d_lt_aswk_reg_4_ ( .D(lt_aswk[4]), .C(clk), .Q(d_lt_aswk[4]) );
  DFFQX1 d_lt_aswk_reg_3_ ( .D(lt_aswk[3]), .C(clk), .Q(d_lt_aswk[3]) );
  DFFQX1 d_lt_aswk_reg_2_ ( .D(lt_aswk[2]), .C(clk), .Q(d_lt_aswk[2]) );
  DFFQX1 d_lt_aswk_reg_1_ ( .D(lt_aswk[1]), .C(clk), .Q(d_lt_aswk[1]) );
  DFFQX1 d_lt_aswk_reg_0_ ( .D(lt_aswk[0]), .C(clk), .Q(d_lt_aswk[0]) );
  DFFQX1 d_lt_gpi_reg_2_ ( .D(lt_gpi[2]), .C(net8975), .Q(d_lt_gpi[2]) );
  DFFQX1 d_regx_addr_reg_4_ ( .D(regx_addr[4]), .C(clk), .Q(d_regx_addr[4]) );
  DFFQX1 d_regx_addr_reg_3_ ( .D(n37), .C(clk), .Q(d_regx_addr[3]) );
  DFFQX1 d_lt_gpi_reg_3_ ( .D(lt_gpi[3]), .C(net8975), .Q(d_lt_gpi[3]) );
  DFFQX1 d_regx_addr_reg_1_ ( .D(regx_addr[1]), .C(clk), .Q(d_regx_addr[1]) );
  DFFQX1 d_regx_addr_reg_6_ ( .D(regx_addr[6]), .C(clk), .Q(d_regx_addr[6]) );
  DFFQX1 d_regx_addr_reg_0_ ( .D(regx_addr[0]), .C(clk), .Q(d_regx_addr[0]) );
  DFFQX1 d_regx_addr_reg_5_ ( .D(regx_addr[5]), .C(clk), .Q(d_regx_addr[5]) );
  DFFRQX1 lt_aswk_reg_5_ ( .D(1'b1), .C(aswclk), .XR(n107), .Q(lt_aswk[5]) );
  DFFRQX1 lt_aswk_reg_4_ ( .D(di_aswk[4]), .C(aswclk), .XR(n107), .Q(
        lt_aswk[4]) );
  DFFRQX1 lt_aswk_reg_3_ ( .D(di_aswk[3]), .C(aswclk), .XR(n107), .Q(
        lt_aswk[3]) );
  DFFRQX1 lt_aswk_reg_2_ ( .D(di_aswk[2]), .C(aswclk), .XR(n107), .Q(
        lt_aswk[2]) );
  DFFRQX1 lt_aswk_reg_1_ ( .D(di_aswk[1]), .C(aswclk), .XR(n107), .Q(
        lt_aswk[1]) );
  DFFRQX1 lt_aswk_reg_0_ ( .D(di_aswk[0]), .C(aswclk), .XR(n107), .Q(
        lt_aswk[0]) );
  DFFRQX1 lt_drp_reg ( .D(di_drposc), .C(detclk), .XR(n52), .Q(lt_drp) );
  AND2XL U3 ( .A(n86), .B(n32), .Y(regx_wrdac[5]) );
  AND2X2 U5 ( .A(n31), .B(n32), .Y(regx_wrdac[8]) );
  OR2X2 U6 ( .A(regx_addr[4]), .B(n33), .Y(n2) );
  AND2XL U7 ( .A(regx_addr[1]), .B(n64), .Y(n31) );
  INVX1 U8 ( .A(n66), .Y(n86) );
  NAND21XL U9 ( .B(regx_addr[1]), .A(n64), .Y(n65) );
  INVX1 U10 ( .A(n91), .Y(n92) );
  NAND21X1 U11 ( .B(n90), .A(n29), .Y(n91) );
  NAND32X1 U12 ( .B(n97), .C(n33), .A(n83), .Y(n94) );
  INVX1 U13 ( .A(regx_addr[6]), .Y(n83) );
  INVX1 U14 ( .A(n85), .Y(n89) );
  NAND21X1 U15 ( .B(n97), .A(n32), .Y(n85) );
  AND2X1 U16 ( .A(n89), .B(n88), .Y(regx_wrdac[7]) );
  AND2X1 U17 ( .A(n92), .B(n102), .Y(regx_wrdac[10]) );
  INVX1 U18 ( .A(n75), .Y(n100) );
  AND2X1 U19 ( .A(n89), .B(n95), .Y(regx_wrdac[4]) );
  AND2X1 U20 ( .A(n89), .B(n104), .Y(regx_wrdac[3]) );
  AND2X1 U21 ( .A(n89), .B(n102), .Y(regx_wrdac[2]) );
  INVX1 U22 ( .A(regx_addr[2]), .Y(n74) );
  INVX1 U23 ( .A(regx_addr[1]), .Y(n73) );
  INVX1 U24 ( .A(regx_addr[5]), .Y(n33) );
  INVX1 U25 ( .A(regx_addr[4]), .Y(n93) );
  INVX1 U26 ( .A(regx_wdat[3]), .Y(n3) );
  INVX1 U27 ( .A(n3), .Y(n4) );
  INVX1 U28 ( .A(n3), .Y(n5) );
  INVX1 U29 ( .A(regx_wdat[6]), .Y(n6) );
  INVX1 U30 ( .A(n6), .Y(n7) );
  INVX1 U31 ( .A(n6), .Y(n8) );
  INVX1 U32 ( .A(regx_wdat[1]), .Y(n9) );
  INVX1 U33 ( .A(n9), .Y(n10) );
  INVX1 U34 ( .A(regx_wdat[4]), .Y(n11) );
  INVX1 U35 ( .A(n11), .Y(n12) );
  INVX1 U36 ( .A(n11), .Y(n13) );
  INVX1 U37 ( .A(regx_wdat[5]), .Y(n14) );
  INVX1 U38 ( .A(n14), .Y(n15) );
  INVX1 U39 ( .A(n14), .Y(n16) );
  INVX1 U40 ( .A(regx_wdat[7]), .Y(n17) );
  INVX1 U41 ( .A(n17), .Y(n18) );
  INVX1 U42 ( .A(n17), .Y(n19) );
  INVX1 U43 ( .A(regx_wdat[2]), .Y(n20) );
  INVX1 U44 ( .A(n20), .Y(n21) );
  INVX1 U45 ( .A(n20), .Y(n22) );
  INVX1 U46 ( .A(regx_wdat[0]), .Y(n23) );
  INVX1 U47 ( .A(n23), .Y(n24) );
  INVXL U48 ( .A(n1048), .Y(n25) );
  INVXL U49 ( .A(n25), .Y(n26) );
  INVX1 U50 ( .A(n109), .Y(n27) );
  INVX1 U51 ( .A(n27), .Y(r_i2crout[5]) );
  BUFX3 U52 ( .A(r_imp_osc), .Y(r_xana[22]) );
  AND2XL U53 ( .A(n92), .B(n104), .Y(regx_wrdac[11]) );
  NOR3X1 U54 ( .A(n37), .B(n94), .C(regx_addr[4]), .Y(n30) );
  AND2XL U55 ( .A(n30), .B(n104), .Y(regx_wrdac[13]) );
  NOR21X4 U56 ( .B(regx_addr[4]), .A(n94), .Y(n29) );
  AND2XL U57 ( .A(n30), .B(n102), .Y(regx_wrdac[12]) );
  NAND32X1 U58 ( .B(regx_addr[0]), .C(n73), .A(n74), .Y(n78) );
  NAND32XL U59 ( .B(regx_addr[1]), .C(n68), .A(n74), .Y(n84) );
  NOR3X2 U60 ( .A(regx_addr[6]), .B(n90), .C(n2), .Y(n32) );
  INVX2 U61 ( .A(regx_addr[3]), .Y(n90) );
  AND2XL U62 ( .A(n96), .B(n104), .Y(regx_wrcvc[1]) );
  AND2XL U63 ( .A(n96), .B(n95), .Y(regx_wrcvc[2]) );
  AND2XL U64 ( .A(n71), .B(n95), .Y(we[26]) );
  AND3XL U65 ( .A(n29), .B(n104), .C(n90), .Y(regx_wrdac[1]) );
  NAND32XL U66 ( .B(n74), .C(n68), .A(n73), .Y(n76) );
  NAND32XL U67 ( .B(n93), .C(n98), .A(n90), .Y(n106) );
  NAND32XL U68 ( .B(n93), .C(n90), .A(n108), .Y(n61) );
  AND2XL U69 ( .A(n86), .B(n103), .Y(we_19) );
  AND2XL U70 ( .A(n67), .B(n86), .Y(we[27]) );
  INVX2 U71 ( .A(regx_addr[0]), .Y(n68) );
  INVX2 U72 ( .A(n70), .Y(n102) );
  INVX1 U73 ( .A(n58), .Y(n55) );
  INVX1 U74 ( .A(n58), .Y(n57) );
  INVX1 U75 ( .A(n59), .Y(n56) );
  INVX1 U76 ( .A(n58), .Y(n48) );
  INVX1 U77 ( .A(n59), .Y(n47) );
  INVX1 U78 ( .A(n58), .Y(n49) );
  INVX1 U79 ( .A(n59), .Y(n46) );
  INVX1 U80 ( .A(n59), .Y(n45) );
  INVX1 U81 ( .A(n58), .Y(n44) );
  INVX1 U82 ( .A(n59), .Y(n43) );
  INVX1 U83 ( .A(n60), .Y(n42) );
  INVX1 U84 ( .A(n58), .Y(n41) );
  INVX1 U85 ( .A(n59), .Y(n40) );
  INVX1 U86 ( .A(n58), .Y(n39) );
  INVX1 U87 ( .A(n60), .Y(n38) );
  INVX1 U88 ( .A(n58), .Y(n50) );
  INVX1 U89 ( .A(n58), .Y(n51) );
  INVX1 U90 ( .A(n59), .Y(n53) );
  INVX1 U91 ( .A(n58), .Y(n52) );
  INVX1 U92 ( .A(n59), .Y(n54) );
  AND2X1 U93 ( .A(n71), .B(n88), .Y(we[29]) );
  INVX1 U94 ( .A(rrstz), .Y(n60) );
  INVX1 U95 ( .A(rrstz), .Y(n58) );
  INVX1 U96 ( .A(rrstz), .Y(n59) );
  INVX1 U97 ( .A(n76), .Y(n88) );
  INVX1 U98 ( .A(n106), .Y(n103) );
  INVX1 U99 ( .A(n72), .Y(n77) );
  NAND21X1 U100 ( .B(n97), .A(n103), .Y(n72) );
  NAND32X1 U101 ( .B(n76), .C(n97), .A(n103), .Y(n1048) );
  INVX1 U102 ( .A(n63), .Y(n71) );
  NAND21X1 U103 ( .B(n97), .A(n67), .Y(n63) );
  AND2XL U104 ( .A(n96), .B(n88), .Y(we_5) );
  AND2X1 U105 ( .A(n67), .B(n31), .Y(we[30]) );
  INVX1 U106 ( .A(n62), .Y(n64) );
  NAND32X1 U107 ( .B(n74), .C(n97), .A(n68), .Y(n62) );
  INVX1 U108 ( .A(n84), .Y(n104) );
  INVX1 U109 ( .A(n78), .Y(n95) );
  AND2X1 U110 ( .A(n102), .B(n103), .Y(regx_hitbst[0]) );
  INVX1 U111 ( .A(n108), .Y(n98) );
  INVX1 U112 ( .A(n79), .Y(we_twlb) );
  NAND21X1 U113 ( .B(n78), .A(n77), .Y(n79) );
  INVX1 U114 ( .A(n81), .Y(n96) );
  NAND21X1 U115 ( .B(n97), .A(n82), .Y(n81) );
  AND2XL U116 ( .A(n101), .B(n104), .Y(regx_wrpwm[1]) );
  AND2X1 U117 ( .A(n101), .B(n102), .Y(regx_wrpwm[0]) );
  AND2X1 U118 ( .A(n96), .B(n102), .Y(regx_wrcvc[0]) );
  INVX1 U119 ( .A(n69), .Y(we[25]) );
  NAND21X1 U120 ( .B(n84), .A(n71), .Y(n69) );
  INVX1 U121 ( .A(n61), .Y(n67) );
  AND2XL U122 ( .A(n104), .B(n103), .Y(regx_hitbst[1]) );
  AND2X1 U123 ( .A(n100), .B(n101), .Y(regx_wrcvc[3]) );
  AND2X1 U124 ( .A(n71), .B(n102), .Y(we[24]) );
  AND2X1 U125 ( .A(n77), .B(n100), .Y(we[23]) );
  AND2X1 U126 ( .A(n96), .B(n100), .Y(we_7) );
  INVX1 U127 ( .A(regx_w), .Y(n97) );
  NAND32XL U128 ( .B(regx_addr[1]), .C(regx_addr[0]), .A(n74), .Y(n70) );
  NAND43X1 U129 ( .B(regx_addr[2]), .C(n68), .D(n97), .A(regx_addr[1]), .Y(n66) );
  NAND32XL U130 ( .B(n74), .C(n73), .A(regx_addr[0]), .Y(n75) );
  NOR2XL U131 ( .A(regx_addr[5]), .B(regx_addr[6]), .Y(n108) );
  INVX1 U132 ( .A(n99), .Y(n101) );
  INVX1 U133 ( .A(n80), .Y(n82) );
  NAND43XL U134 ( .B(regx_addr[5]), .C(regx_addr[6]), .D(n37), .A(n93), .Y(n80) );
  OAI31XL U135 ( .A(n17), .B(n8), .C(n26), .D(n1049), .Y(i2c_mode_upd) );
  OAI21X1 U136 ( .B(n1050), .C(n1051), .A(bus_idle), .Y(n1049) );
  NAND3X1 U137 ( .A(n1052), .B(n1053), .C(n1054), .Y(n1051) );
  NOR4XL U138 ( .A(n1058), .B(n1059), .C(regx_wdat[3]), .D(n21), .Y(N8) );
  NAND3X1 U139 ( .A(n14), .B(n9), .C(n11), .Y(n1059) );
  NAND43X1 U140 ( .B(n106), .C(n6), .D(regx_addr[0]), .A(n105), .Y(n1058) );
  AND2X1 U141 ( .A(regx_w), .B(regx_wdat[0]), .Y(n1060) );
  BUFX3 U142 ( .A(n24), .Y(wd_twlb[0]) );
  BUFX3 U143 ( .A(n10), .Y(wd_twlb[1]) );
  ENOX1 U144 ( .A(n1048), .B(n9), .C(n26), .D(lt_reg15_5_0[1]), .Y(
        i2c_mode_wdat[1]) );
  ENOX1 U145 ( .A(n26), .B(n11), .C(n1048), .D(lt_reg15_5_0[4]), .Y(
        i2c_mode_wdat[4]) );
  ENOX1 U146 ( .A(n1048), .B(n14), .C(n26), .D(lt_reg15_5_0[5]), .Y(
        i2c_mode_wdat[5]) );
  NAND4X1 U147 ( .A(n1055), .B(n1056), .C(n1057), .D(n26), .Y(n1050) );
  XNOR2XL U148 ( .A(r_i2crout[3]), .B(lt_reg15_5_0[3]), .Y(n1055) );
  XNOR2XL U149 ( .A(r_i2crout[4]), .B(lt_reg15_5_0[4]), .Y(n1056) );
  XNOR2XL U150 ( .A(n109), .B(lt_reg15_5_0[5]), .Y(n1057) );
  AO22X1 U151 ( .A(n25), .B(n24), .C(n1048), .D(lt_reg15_5_0[0]), .Y(
        i2c_mode_wdat[0]) );
  AO22X1 U152 ( .A(n25), .B(n22), .C(n26), .D(lt_reg15_5_0[2]), .Y(
        i2c_mode_wdat[2]) );
  AO22X1 U153 ( .A(n25), .B(n4), .C(n1048), .D(lt_reg15_5_0[3]), .Y(
        i2c_mode_wdat[3]) );
  XNOR2XL U154 ( .A(reg1E[3]), .B(n1047), .Y(r_xana[19]) );
  XNOR2XL U155 ( .A(reg1E[2]), .B(n1047), .Y(r_xana[18]) );
  NAND2X1 U156 ( .A(r_xana[20]), .B(di_drposc), .Y(n1047) );
  XNOR2XL U157 ( .A(r_i2crout[2]), .B(lt_reg15_5_0[2]), .Y(n1052) );
  XNOR2XL U158 ( .A(r_i2crout[0]), .B(lt_reg15_5_0[0]), .Y(n1053) );
  XNOR2XL U159 ( .A(r_i2crout[1]), .B(lt_reg15_5_0[1]), .Y(n1054) );
  INVX1 U160 ( .A(n1061), .Y(n107) );
  OAI21BX1 U161 ( .C(d_we16), .B(atpg_en), .A(n53), .Y(n1061) );
  AND2X2 U162 ( .A(n89), .B(n100), .Y(regx_wrdac[9]) );
  BUFXL U163 ( .A(regx_addr[3]), .Y(n37) );
  AND3X1 U164 ( .A(n29), .B(n102), .C(n90), .Y(regx_wrdac[0]) );
  NAND43XL U165 ( .B(regx_addr[4]), .C(n98), .D(n97), .A(n37), .Y(n99) );
  AND2XL U166 ( .A(n67), .B(n87), .Y(we[28]) );
  AND2XL U167 ( .A(n87), .B(n82), .Y(we_4) );
  AND2X2 U168 ( .A(n87), .B(n32), .Y(regx_wrdac[6]) );
  INVX3 U169 ( .A(n65), .Y(n87) );
  AND4XL U170 ( .A(n1060), .B(regx_addr[2]), .C(n18), .D(regx_addr[1]), .Y(
        n105) );
endmodule


module regx_a0_DW_rightsh_0 ( A, DATA_TC, SH, B );
  input [1023:0] A;
  input [9:0] SH;
  output [1023:0] B;
  input DATA_TC;
  wire   n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171,
         n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181,
         n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191,
         n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201,
         n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211,
         n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221,
         n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231,
         n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241,
         n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251,
         n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261,
         n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271,
         n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281,
         n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291,
         n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301,
         n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311,
         n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321,
         n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331,
         n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341,
         n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351,
         n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361,
         n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371,
         n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381,
         n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391,
         n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401,
         n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411,
         n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421,
         n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431,
         n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441,
         n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451,
         n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461,
         n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471,
         n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481,
         n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491,
         n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501,
         n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511,
         n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521,
         n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531,
         n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541,
         n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551,
         n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561,
         n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571,
         n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581,
         n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591,
         n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601,
         n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611,
         n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621,
         n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631,
         n3632;

  BUFX3 U2125 ( .A(SH[6]), .Y(n3162) );
  BUFX3 U2126 ( .A(SH[5]), .Y(n3163) );
  INVX1 U2127 ( .A(n3197), .Y(n3184) );
  INVX1 U2128 ( .A(n3196), .Y(n3186) );
  INVX1 U2129 ( .A(n3197), .Y(n3185) );
  INVX1 U2130 ( .A(n3194), .Y(n3193) );
  INVX1 U2131 ( .A(n3197), .Y(n3183) );
  INVX1 U2132 ( .A(n3198), .Y(n3181) );
  INVX1 U2133 ( .A(n3198), .Y(n3180) );
  INVX1 U2134 ( .A(n3198), .Y(n3182) );
  INVX1 U2135 ( .A(n3238), .Y(n3213) );
  INVX1 U2136 ( .A(n3238), .Y(n3214) );
  INVX1 U2137 ( .A(n3196), .Y(n3187) );
  INVX1 U2138 ( .A(n3233), .Y(n3222) );
  INVX1 U2139 ( .A(n3234), .Y(n3220) );
  INVX1 U2140 ( .A(n3233), .Y(n3223) );
  INVX1 U2141 ( .A(n3238), .Y(n3221) );
  INVX1 U2142 ( .A(n3233), .Y(n3215) );
  INVX1 U2143 ( .A(n3234), .Y(n3225) );
  INVX1 U2144 ( .A(n3234), .Y(n3226) );
  INVX1 U2145 ( .A(n3196), .Y(n3188) );
  INVX1 U2146 ( .A(n3234), .Y(n3231) );
  INVX1 U2147 ( .A(n3234), .Y(n3230) );
  INVX1 U2148 ( .A(n3233), .Y(n3229) );
  INVX1 U2149 ( .A(n3195), .Y(n3189) );
  INVX1 U2150 ( .A(n3234), .Y(n3224) );
  INVX1 U2151 ( .A(n3232), .Y(n3219) );
  INVX1 U2152 ( .A(n3232), .Y(n3217) );
  INVX1 U2153 ( .A(n3234), .Y(n3216) );
  INVX1 U2154 ( .A(n3232), .Y(n3218) );
  INVX1 U2155 ( .A(n3238), .Y(n3227) );
  INVX1 U2156 ( .A(n3238), .Y(n3228) );
  INVX1 U2157 ( .A(n3198), .Y(n3192) );
  INVX1 U2158 ( .A(n3198), .Y(n3191) );
  INVX1 U2159 ( .A(n3198), .Y(n3190) );
  INVX1 U2160 ( .A(n3208), .Y(n3197) );
  INVX1 U2161 ( .A(n3209), .Y(n3194) );
  INVX1 U2162 ( .A(n3208), .Y(n3196) );
  INVX1 U2163 ( .A(n3237), .Y(n3232) );
  INVX1 U2164 ( .A(n3208), .Y(n3198) );
  INVX1 U2165 ( .A(n3236), .Y(n3233) );
  INVX1 U2166 ( .A(n3235), .Y(n3234) );
  INVX1 U2167 ( .A(n3209), .Y(n3195) );
  INVX1 U2168 ( .A(n3207), .Y(n3199) );
  INVX1 U2169 ( .A(n3206), .Y(n3201) );
  INVX1 U2170 ( .A(n3207), .Y(n3200) );
  INVX1 U2171 ( .A(n3205), .Y(n3202) );
  INVX1 U2172 ( .A(n3210), .Y(n3208) );
  INVX1 U2173 ( .A(n3210), .Y(n3209) );
  INVX1 U2174 ( .A(n3171), .Y(n3170) );
  INVX1 U2175 ( .A(n3210), .Y(n3207) );
  INVX1 U2176 ( .A(n3211), .Y(n3206) );
  INVX1 U2177 ( .A(n3238), .Y(n3235) );
  INVX1 U2178 ( .A(n3238), .Y(n3236) );
  INVX1 U2179 ( .A(n3238), .Y(n3237) );
  INVX1 U2180 ( .A(n3205), .Y(n3203) );
  INVX1 U2181 ( .A(n3205), .Y(n3204) );
  INVX1 U2182 ( .A(n3171), .Y(n3164) );
  INVX1 U2183 ( .A(n3171), .Y(n3165) );
  INVX1 U2184 ( .A(n3171), .Y(n3167) );
  INVX1 U2185 ( .A(n3171), .Y(n3168) );
  INVX1 U2186 ( .A(n3179), .Y(n3177) );
  INVX1 U2187 ( .A(n3179), .Y(n3178) );
  INVX1 U2188 ( .A(n3172), .Y(n3169) );
  INVX1 U2189 ( .A(n3179), .Y(n3174) );
  INVX1 U2190 ( .A(n3179), .Y(n3175) );
  INVX1 U2191 ( .A(n3179), .Y(n3176) );
  INVX1 U2192 ( .A(n3171), .Y(n3166) );
  INVX1 U2193 ( .A(SH[8]), .Y(n3210) );
  INVX1 U2194 ( .A(n3212), .Y(n3205) );
  INVX1 U2195 ( .A(SH[8]), .Y(n3212) );
  INVX1 U2196 ( .A(SH[8]), .Y(n3211) );
  INVX1 U2197 ( .A(SH[9]), .Y(n3238) );
  INVX1 U2198 ( .A(n3179), .Y(n3173) );
  INVX1 U2199 ( .A(SH[4]), .Y(n3179) );
  INVX1 U2200 ( .A(SH[3]), .Y(n3171) );
  INVX1 U2201 ( .A(SH[3]), .Y(n3172) );
  MUX2IX1 U2202 ( .D0(n3239), .D1(n3240), .S(SH[7]), .Y(B[7]) );
  MUX4X1 U2203 ( .D0(n3241), .D1(n3242), .D2(n3243), .D3(n3244), .S0(SH[5]), 
        .S1(SH[6]), .Y(n3240) );
  MUX4X1 U2204 ( .D0(n3245), .D1(n3246), .D2(n3247), .D3(n3248), .S0(n3173), 
        .S1(n3167), .Y(n3244) );
  NOR3XL U2205 ( .A(A[255]), .B(n3215), .C(n3189), .Y(n3248) );
  NOR3XL U2206 ( .A(A[239]), .B(n3223), .C(n3189), .Y(n3247) );
  NOR3XL U2207 ( .A(A[247]), .B(n3220), .C(n3193), .Y(n3246) );
  NOR3XL U2208 ( .A(A[231]), .B(n3220), .C(n3193), .Y(n3245) );
  MUX4X1 U2209 ( .D0(n3249), .D1(n3250), .D2(n3251), .D3(n3252), .S0(n3173), 
        .S1(n3169), .Y(n3243) );
  NOR3XL U2210 ( .A(A[223]), .B(n3221), .C(n3193), .Y(n3252) );
  AOI21X1 U2211 ( .B(A[207]), .C(n3199), .A(n3213), .Y(n3251) );
  AOI21X1 U2212 ( .B(A[215]), .C(n3199), .A(n3213), .Y(n3250) );
  AOI21X1 U2213 ( .B(A[199]), .C(n3199), .A(n3213), .Y(n3249) );
  MUX3X1 U2214 ( .D0(n3253), .D1(n3254), .D2(n3255), .S0(n3169), .S1(SH[4]), 
        .Y(n3242) );
  AOI211X1 U2215 ( .C(n3170), .D(A[191]), .A(n3214), .B(n3187), .Y(n3255) );
  NOR3XL U2216 ( .A(A[175]), .B(n3221), .C(n3193), .Y(n3254) );
  NOR3XL U2217 ( .A(A[167]), .B(n3221), .C(n3193), .Y(n3253) );
  MUX4X1 U2218 ( .D0(n3256), .D1(n3257), .D2(n3258), .D3(n3259), .S0(n3173), 
        .S1(n3168), .Y(n3241) );
  NOR3XL U2219 ( .A(A[159]), .B(n3221), .C(n3193), .Y(n3259) );
  NOR21XL U2220 ( .B(n3260), .A(n3231), .Y(n3258) );
  MUX2IX1 U2221 ( .D0(A[143]), .D1(A[399]), .S(n3185), .Y(n3260) );
  NOR21XL U2222 ( .B(n3261), .A(n3230), .Y(n3257) );
  MUX2IX1 U2223 ( .D0(A[151]), .D1(A[407]), .S(n3184), .Y(n3261) );
  NOR21XL U2224 ( .B(n3262), .A(n3230), .Y(n3256) );
  MUX2IX1 U2225 ( .D0(A[135]), .D1(A[391]), .S(n3186), .Y(n3262) );
  MUX4X1 U2226 ( .D0(n3263), .D1(n3264), .D2(n3265), .D3(n3266), .S0(SH[6]), 
        .S1(SH[5]), .Y(n3239) );
  MUX4X1 U2227 ( .D0(n3267), .D1(n3268), .D2(n3269), .D3(n3270), .S0(n3173), 
        .S1(n3168), .Y(n3266) );
  NOR21XL U2228 ( .B(n3271), .A(n3230), .Y(n3270) );
  MUX2IX1 U2229 ( .D0(A[127]), .D1(A[383]), .S(n3185), .Y(n3271) );
  NOR3XL U2230 ( .A(n3201), .B(n3221), .C(A[367]), .Y(n3269) );
  NOR3XL U2231 ( .A(n3204), .B(n3221), .C(A[375]), .Y(n3268) );
  NOR3XL U2232 ( .A(n3204), .B(n3221), .C(A[359]), .Y(n3267) );
  MUX3X1 U2233 ( .D0(n3272), .D1(n3273), .D2(n3274), .S0(n3169), .S1(SH[4]), 
        .Y(n3265) );
  NOR4XL U2234 ( .A(n3226), .B(n3188), .C(A[63]), .D(n3172), .Y(n3274) );
  NOR3XL U2235 ( .A(A[47]), .B(n3221), .C(n3193), .Y(n3273) );
  NOR3XL U2236 ( .A(A[39]), .B(n3221), .C(n3193), .Y(n3272) );
  MUX4X1 U2237 ( .D0(n3275), .D1(n3276), .D2(n3277), .D3(n3278), .S0(n3164), 
        .S1(n3177), .Y(n3264) );
  NOR3XL U2238 ( .A(n3203), .B(n3221), .C(A[351]), .Y(n3278) );
  NOR3XL U2239 ( .A(n3203), .B(n3222), .C(A[343]), .Y(n3277) );
  NOR21XL U2240 ( .B(n3279), .A(n3229), .Y(n3276) );
  MUX2IX1 U2241 ( .D0(A[79]), .D1(A[335]), .S(n3185), .Y(n3279) );
  NOR21XL U2242 ( .B(n3280), .A(n3229), .Y(n3275) );
  MUX2IX1 U2243 ( .D0(A[71]), .D1(A[327]), .S(n3186), .Y(n3280) );
  MUX2X1 U2244 ( .D0(n3281), .D1(n3282), .S(n3178), .Y(n3263) );
  NOR4XL U2245 ( .A(n3225), .B(n3187), .C(n3170), .D(A[23]), .Y(n3282) );
  MUX2IX1 U2246 ( .D0(n3283), .D1(n3284), .S(n3165), .Y(n3281) );
  NAND2X1 U2247 ( .A(n3285), .B(n3238), .Y(n3284) );
  MUX2IX1 U2248 ( .D0(A[15]), .D1(A[271]), .S(n3186), .Y(n3285) );
  NAND2X1 U2249 ( .A(n3286), .B(n3232), .Y(n3283) );
  MUX2IX1 U2250 ( .D0(A[7]), .D1(A[263]), .S(n3186), .Y(n3286) );
  MUX2IX1 U2251 ( .D0(n3287), .D1(n3288), .S(SH[7]), .Y(B[6]) );
  MUX4X1 U2252 ( .D0(n3289), .D1(n3290), .D2(n3291), .D3(n3292), .S0(SH[5]), 
        .S1(n3162), .Y(n3288) );
  MUX4X1 U2253 ( .D0(n3293), .D1(n3294), .D2(n3295), .D3(n3296), .S0(n3173), 
        .S1(n3166), .Y(n3292) );
  NOR3XL U2254 ( .A(A[254]), .B(n3222), .C(n3206), .Y(n3296) );
  NOR3XL U2255 ( .A(A[238]), .B(n3222), .C(n3205), .Y(n3295) );
  NOR3XL U2256 ( .A(A[246]), .B(n3222), .C(n3207), .Y(n3294) );
  NOR3XL U2257 ( .A(A[230]), .B(n3222), .C(n3207), .Y(n3293) );
  MUX4X1 U2258 ( .D0(n3297), .D1(n3298), .D2(n3299), .D3(n3300), .S0(n3173), 
        .S1(n3166), .Y(n3291) );
  NOR3XL U2259 ( .A(A[222]), .B(n3222), .C(n3207), .Y(n3300) );
  AOI21X1 U2260 ( .B(A[206]), .C(n3202), .A(n3213), .Y(n3299) );
  AOI21X1 U2261 ( .B(A[214]), .C(n3211), .A(n3213), .Y(n3298) );
  AOI21X1 U2262 ( .B(A[198]), .C(n3200), .A(n3214), .Y(n3297) );
  MUX2X1 U2263 ( .D0(n3301), .D1(n3302), .S(n3178), .Y(n3290) );
  AOI211X1 U2264 ( .C(n3170), .D(A[190]), .A(SH[9]), .B(n3187), .Y(n3302) );
  AOI211X1 U2265 ( .C(A[166]), .D(n3171), .A(SH[9]), .B(n3187), .Y(n3301) );
  MUX4X1 U2266 ( .D0(n3303), .D1(n3304), .D2(n3305), .D3(n3306), .S0(n3174), 
        .S1(n3165), .Y(n3289) );
  NOR3XL U2267 ( .A(A[158]), .B(n3222), .C(n3205), .Y(n3306) );
  NOR21XL U2268 ( .B(n3307), .A(n3228), .Y(n3305) );
  MUX2IX1 U2269 ( .D0(A[142]), .D1(A[398]), .S(n3185), .Y(n3307) );
  NOR21XL U2270 ( .B(n3308), .A(n3228), .Y(n3304) );
  MUX2IX1 U2271 ( .D0(A[150]), .D1(A[406]), .S(n3186), .Y(n3308) );
  NOR21XL U2272 ( .B(n3309), .A(n3229), .Y(n3303) );
  MUX2IX1 U2273 ( .D0(A[134]), .D1(A[390]), .S(n3184), .Y(n3309) );
  MUX4X1 U2274 ( .D0(n3310), .D1(n3311), .D2(n3312), .D3(n3313), .S0(SH[6]), 
        .S1(n3163), .Y(n3287) );
  MUX4X1 U2275 ( .D0(n3314), .D1(n3315), .D2(n3316), .D3(n3317), .S0(n3174), 
        .S1(n3165), .Y(n3313) );
  NOR21XL U2276 ( .B(n3318), .A(n3227), .Y(n3317) );
  MUX2IX1 U2277 ( .D0(A[126]), .D1(A[382]), .S(n3185), .Y(n3318) );
  NOR3XL U2278 ( .A(n3203), .B(n3222), .C(A[366]), .Y(n3316) );
  NOR3XL U2279 ( .A(n3203), .B(n3222), .C(A[374]), .Y(n3315) );
  NOR3XL U2280 ( .A(n3211), .B(n3222), .C(A[358]), .Y(n3314) );
  MUX3X1 U2281 ( .D0(n3319), .D1(n3320), .D2(n3321), .S0(n3169), .S1(n3178), 
        .Y(n3312) );
  NOR4XL U2282 ( .A(n3225), .B(n3187), .C(A[62]), .D(n3172), .Y(n3321) );
  NOR3XL U2283 ( .A(A[46]), .B(n3235), .C(n3207), .Y(n3320) );
  NOR3XL U2284 ( .A(A[38]), .B(n3237), .C(n3207), .Y(n3319) );
  MUX4X1 U2285 ( .D0(n3322), .D1(n3323), .D2(n3324), .D3(n3325), .S0(n3164), 
        .S1(n3176), .Y(n3311) );
  NOR3XL U2286 ( .A(n3202), .B(n3235), .C(A[350]), .Y(n3325) );
  NOR3XL U2287 ( .A(n3204), .B(n3235), .C(A[342]), .Y(n3324) );
  NOR21XL U2288 ( .B(n3326), .A(n3228), .Y(n3323) );
  MUX2IX1 U2289 ( .D0(A[78]), .D1(A[334]), .S(n3184), .Y(n3326) );
  NOR21XL U2290 ( .B(n3327), .A(n3227), .Y(n3322) );
  MUX2IX1 U2291 ( .D0(A[70]), .D1(A[326]), .S(n3185), .Y(n3327) );
  MUX2X1 U2292 ( .D0(n3328), .D1(n3329), .S(n3178), .Y(n3310) );
  NOR4XL U2293 ( .A(n3225), .B(n3187), .C(SH[3]), .D(A[22]), .Y(n3329) );
  MUX2IX1 U2294 ( .D0(n3330), .D1(n3331), .S(n3165), .Y(n3328) );
  NAND2X1 U2295 ( .A(n3332), .B(n3232), .Y(n3331) );
  MUX2IX1 U2296 ( .D0(A[14]), .D1(A[270]), .S(n3185), .Y(n3332) );
  NAND2X1 U2297 ( .A(n3333), .B(n3232), .Y(n3330) );
  MUX2IX1 U2298 ( .D0(A[6]), .D1(A[262]), .S(n3185), .Y(n3333) );
  MUX2IX1 U2299 ( .D0(n3334), .D1(n3335), .S(SH[7]), .Y(B[5]) );
  MUX4X1 U2300 ( .D0(n3336), .D1(n3337), .D2(n3338), .D3(n3339), .S0(SH[5]), 
        .S1(n3162), .Y(n3335) );
  MUX3X1 U2301 ( .D0(n3340), .D1(n3341), .D2(n3342), .S0(n3169), .S1(n3178), 
        .Y(n3339) );
  AOI211X1 U2302 ( .C(A[245]), .D(n3172), .A(n3214), .B(n3187), .Y(n3342) );
  NOR3XL U2303 ( .A(A[237]), .B(n3237), .C(n3205), .Y(n3341) );
  NOR3XL U2304 ( .A(A[229]), .B(n3237), .C(n3207), .Y(n3340) );
  MUX4X1 U2305 ( .D0(n3343), .D1(n3344), .D2(n3345), .D3(n3346), .S0(n3174), 
        .S1(n3166), .Y(n3338) );
  NOR3XL U2306 ( .A(A[221]), .B(n3237), .C(n3206), .Y(n3346) );
  AOI21X1 U2307 ( .B(A[205]), .C(n3200), .A(n3213), .Y(n3345) );
  AOI21X1 U2308 ( .B(A[213]), .C(n3200), .A(n3213), .Y(n3344) );
  AOI21X1 U2309 ( .B(A[197]), .C(n3200), .A(n3214), .Y(n3343) );
  MUX4X1 U2310 ( .D0(n3347), .D1(n3348), .D2(n3349), .D3(n3350), .S0(n3174), 
        .S1(n3165), .Y(n3337) );
  NOR3XL U2311 ( .A(A[189]), .B(n3235), .C(n3206), .Y(n3350) );
  NOR3XL U2312 ( .A(A[173]), .B(n3235), .C(n3205), .Y(n3349) );
  NOR3XL U2313 ( .A(A[181]), .B(n3235), .C(n3206), .Y(n3348) );
  NOR3XL U2314 ( .A(A[165]), .B(n3223), .C(n3206), .Y(n3347) );
  MUX4X1 U2315 ( .D0(n3351), .D1(n3352), .D2(n3353), .D3(n3354), .S0(n3174), 
        .S1(n3166), .Y(n3336) );
  NOR3XL U2316 ( .A(A[157]), .B(n3223), .C(n3206), .Y(n3354) );
  NOR21XL U2317 ( .B(n3355), .A(n3228), .Y(n3353) );
  MUX2IX1 U2318 ( .D0(A[141]), .D1(A[397]), .S(n3184), .Y(n3355) );
  NOR21XL U2319 ( .B(n3356), .A(n3226), .Y(n3352) );
  MUX2IX1 U2320 ( .D0(A[149]), .D1(A[405]), .S(n3184), .Y(n3356) );
  NOR21XL U2321 ( .B(n3357), .A(n3226), .Y(n3351) );
  MUX2IX1 U2322 ( .D0(A[133]), .D1(A[389]), .S(n3184), .Y(n3357) );
  MUX4X1 U2323 ( .D0(n3358), .D1(n3359), .D2(n3360), .D3(n3361), .S0(n3162), 
        .S1(n3163), .Y(n3334) );
  MUX4X1 U2324 ( .D0(n3362), .D1(n3363), .D2(n3364), .D3(n3365), .S0(n3174), 
        .S1(n3166), .Y(n3361) );
  NOR21XL U2325 ( .B(n3366), .A(n3226), .Y(n3365) );
  MUX2IX1 U2326 ( .D0(A[125]), .D1(A[381]), .S(n3183), .Y(n3366) );
  NOR3XL U2327 ( .A(n3200), .B(n3223), .C(A[365]), .Y(n3364) );
  NOR3XL U2328 ( .A(n3202), .B(n3223), .C(A[373]), .Y(n3363) );
  NOR3XL U2329 ( .A(n3202), .B(n3223), .C(A[357]), .Y(n3362) );
  MUX3X1 U2330 ( .D0(n3367), .D1(n3368), .D2(n3369), .S0(n3169), .S1(n3178), 
        .Y(n3360) );
  NOR4XL U2331 ( .A(n3225), .B(n3187), .C(A[61]), .D(n3172), .Y(n3369) );
  NOR3XL U2332 ( .A(A[45]), .B(n3223), .C(n3205), .Y(n3368) );
  NOR3XL U2333 ( .A(A[37]), .B(n3223), .C(n3205), .Y(n3367) );
  MUX4X1 U2334 ( .D0(n3370), .D1(n3371), .D2(n3372), .D3(n3373), .S0(n3164), 
        .S1(n3177), .Y(n3359) );
  NOR3XL U2335 ( .A(n3202), .B(n3224), .C(A[349]), .Y(n3373) );
  NOR3XL U2336 ( .A(n3202), .B(n3224), .C(A[341]), .Y(n3372) );
  NOR21XL U2337 ( .B(n3374), .A(n3227), .Y(n3371) );
  MUX2IX1 U2338 ( .D0(A[77]), .D1(A[333]), .S(n3183), .Y(n3374) );
  NOR21XL U2339 ( .B(n3375), .A(n3229), .Y(n3370) );
  MUX2IX1 U2340 ( .D0(A[69]), .D1(A[325]), .S(n3184), .Y(n3375) );
  MUX2X1 U2341 ( .D0(n3376), .D1(n3377), .S(n3178), .Y(n3358) );
  NOR4XL U2342 ( .A(n3226), .B(n3187), .C(n3170), .D(A[21]), .Y(n3377) );
  MUX2IX1 U2343 ( .D0(n3378), .D1(n3379), .S(n3165), .Y(n3376) );
  NAND2X1 U2344 ( .A(n3380), .B(n3233), .Y(n3379) );
  MUX2IX1 U2345 ( .D0(A[13]), .D1(A[269]), .S(n3183), .Y(n3380) );
  NAND2X1 U2346 ( .A(n3381), .B(n3234), .Y(n3378) );
  MUX2IX1 U2347 ( .D0(A[5]), .D1(A[261]), .S(n3183), .Y(n3381) );
  MUX2IX1 U2348 ( .D0(n3382), .D1(n3383), .S(SH[7]), .Y(B[4]) );
  MUX4X1 U2349 ( .D0(n3384), .D1(n3385), .D2(n3386), .D3(n3387), .S0(n3163), 
        .S1(n3162), .Y(n3383) );
  MUX4X1 U2350 ( .D0(n3388), .D1(n3389), .D2(n3390), .D3(n3391), .S0(n3175), 
        .S1(n3165), .Y(n3387) );
  NOR3XL U2351 ( .A(A[252]), .B(n3224), .C(n3205), .Y(n3391) );
  NOR3XL U2352 ( .A(A[236]), .B(n3224), .C(n3206), .Y(n3390) );
  NOR3XL U2353 ( .A(A[244]), .B(n3224), .C(n3192), .Y(n3389) );
  NOR3XL U2354 ( .A(A[228]), .B(n3223), .C(n3192), .Y(n3388) );
  MUX4X1 U2355 ( .D0(n3392), .D1(n3393), .D2(n3394), .D3(n3395), .S0(n3175), 
        .S1(n3166), .Y(n3386) );
  NOR3XL U2356 ( .A(A[220]), .B(n3224), .C(n3192), .Y(n3395) );
  AOI21X1 U2357 ( .B(A[204]), .C(n3200), .A(n3214), .Y(n3394) );
  AOI21X1 U2358 ( .B(A[212]), .C(n3204), .A(n3214), .Y(n3393) );
  AOI21X1 U2359 ( .B(A[196]), .C(n3198), .A(n3214), .Y(n3392) );
  MUX4X1 U2360 ( .D0(n3396), .D1(n3397), .D2(n3398), .D3(n3399), .S0(n3173), 
        .S1(n3166), .Y(n3385) );
  NOR3XL U2361 ( .A(A[188]), .B(n3223), .C(n3192), .Y(n3399) );
  NOR3XL U2362 ( .A(A[172]), .B(n3224), .C(n3192), .Y(n3398) );
  NOR3XL U2363 ( .A(A[180]), .B(n3224), .C(n3192), .Y(n3397) );
  NOR3XL U2364 ( .A(A[164]), .B(n3224), .C(n3192), .Y(n3396) );
  MUX4X1 U2365 ( .D0(n3400), .D1(n3401), .D2(n3402), .D3(n3403), .S0(n3175), 
        .S1(n3166), .Y(n3384) );
  NOR3XL U2366 ( .A(A[156]), .B(n3224), .C(n3192), .Y(n3403) );
  NOR21XL U2367 ( .B(n3404), .A(n3231), .Y(n3402) );
  MUX2IX1 U2368 ( .D0(A[140]), .D1(A[396]), .S(n3182), .Y(n3404) );
  NOR21XL U2369 ( .B(n3405), .A(n3231), .Y(n3401) );
  MUX2IX1 U2370 ( .D0(A[148]), .D1(A[404]), .S(n3182), .Y(n3405) );
  NOR21XL U2371 ( .B(n3406), .A(n3231), .Y(n3400) );
  MUX2IX1 U2372 ( .D0(A[132]), .D1(A[388]), .S(n3182), .Y(n3406) );
  MUX4X1 U2373 ( .D0(n3407), .D1(n3408), .D2(n3409), .D3(n3410), .S0(n3162), 
        .S1(n3163), .Y(n3382) );
  MUX4X1 U2374 ( .D0(n3411), .D1(n3412), .D2(n3413), .D3(n3414), .S0(n3175), 
        .S1(n3166), .Y(n3410) );
  NOR21XL U2375 ( .B(n3415), .A(n3231), .Y(n3414) );
  MUX2IX1 U2376 ( .D0(A[124]), .D1(A[380]), .S(n3182), .Y(n3415) );
  NOR3XL U2377 ( .A(n3212), .B(n3220), .C(A[364]), .Y(n3413) );
  NOR3XL U2378 ( .A(n3204), .B(n3220), .C(A[372]), .Y(n3412) );
  NOR3XL U2379 ( .A(n3204), .B(n3220), .C(A[356]), .Y(n3411) );
  MUX3X1 U2380 ( .D0(n3416), .D1(n3417), .D2(n3418), .S0(n3169), .S1(n3178), 
        .Y(n3409) );
  NOR4XL U2381 ( .A(n3226), .B(n3188), .C(A[60]), .D(n3172), .Y(n3418) );
  NOR3XL U2382 ( .A(A[44]), .B(n3220), .C(n3192), .Y(n3417) );
  NOR3XL U2383 ( .A(A[36]), .B(n3220), .C(n3192), .Y(n3416) );
  MUX4X1 U2384 ( .D0(n3419), .D1(n3420), .D2(n3421), .D3(n3422), .S0(n3164), 
        .S1(n3177), .Y(n3408) );
  NOR3XL U2385 ( .A(n3211), .B(n3220), .C(A[348]), .Y(n3422) );
  NOR3XL U2386 ( .A(n3203), .B(n3220), .C(A[340]), .Y(n3421) );
  NOR21XL U2387 ( .B(n3423), .A(n3230), .Y(n3420) );
  MUX2IX1 U2388 ( .D0(A[76]), .D1(A[332]), .S(n3182), .Y(n3423) );
  NOR21XL U2389 ( .B(n3424), .A(n3230), .Y(n3419) );
  MUX2IX1 U2390 ( .D0(A[68]), .D1(A[324]), .S(n3182), .Y(n3424) );
  MUX2X1 U2391 ( .D0(n3425), .D1(n3426), .S(n3177), .Y(n3407) );
  NOR4XL U2392 ( .A(n3226), .B(n3188), .C(n3170), .D(A[20]), .Y(n3426) );
  MUX2IX1 U2393 ( .D0(n3427), .D1(n3428), .S(n3165), .Y(n3425) );
  NAND2X1 U2394 ( .A(n3429), .B(n3238), .Y(n3428) );
  MUX2IX1 U2395 ( .D0(A[12]), .D1(A[268]), .S(n3182), .Y(n3429) );
  NAND2X1 U2396 ( .A(n3430), .B(n3232), .Y(n3427) );
  MUX2IX1 U2397 ( .D0(A[4]), .D1(A[260]), .S(n3181), .Y(n3430) );
  MUX2IX1 U2398 ( .D0(n3431), .D1(n3432), .S(SH[7]), .Y(B[3]) );
  MUX4X1 U2399 ( .D0(n3433), .D1(n3434), .D2(n3435), .D3(n3436), .S0(SH[5]), 
        .S1(SH[6]), .Y(n3432) );
  MUX4X1 U2400 ( .D0(n3437), .D1(n3438), .D2(n3439), .D3(n3440), .S0(n3175), 
        .S1(n3167), .Y(n3436) );
  NOR3XL U2401 ( .A(A[251]), .B(n3236), .C(n3191), .Y(n3440) );
  NOR3XL U2402 ( .A(A[235]), .B(n3236), .C(n3191), .Y(n3439) );
  NOR3XL U2403 ( .A(A[243]), .B(n3237), .C(n3191), .Y(n3438) );
  NOR3XL U2404 ( .A(A[227]), .B(SH[9]), .C(n3191), .Y(n3437) );
  MUX4X1 U2405 ( .D0(n3441), .D1(n3442), .D2(n3443), .D3(n3444), .S0(n3175), 
        .S1(n3167), .Y(n3435) );
  NOR3XL U2406 ( .A(A[219]), .B(n3236), .C(n3191), .Y(n3444) );
  AOI21X1 U2407 ( .B(A[203]), .C(n3198), .A(n3213), .Y(n3443) );
  AOI21X1 U2408 ( .B(A[211]), .C(n3201), .A(n3214), .Y(n3442) );
  AOI21X1 U2409 ( .B(A[195]), .C(n3200), .A(n3214), .Y(n3441) );
  MUX4X1 U2410 ( .D0(n3445), .D1(n3446), .D2(n3447), .D3(n3448), .S0(n3174), 
        .S1(n3166), .Y(n3434) );
  NOR3XL U2411 ( .A(A[187]), .B(n3237), .C(n3191), .Y(n3448) );
  NOR3XL U2412 ( .A(A[171]), .B(SH[9]), .C(n3191), .Y(n3447) );
  NOR3XL U2413 ( .A(A[179]), .B(n3219), .C(n3191), .Y(n3446) );
  NOR3XL U2414 ( .A(A[163]), .B(n3235), .C(n3191), .Y(n3445) );
  MUX4X1 U2415 ( .D0(n3449), .D1(n3450), .D2(n3451), .D3(n3452), .S0(n3175), 
        .S1(n3167), .Y(n3433) );
  NOR3XL U2416 ( .A(A[155]), .B(n3219), .C(n3191), .Y(n3452) );
  NOR21XL U2417 ( .B(n3453), .A(n3227), .Y(n3451) );
  MUX2IX1 U2418 ( .D0(A[139]), .D1(A[395]), .S(n3181), .Y(n3453) );
  NOR21XL U2419 ( .B(n3454), .A(n3227), .Y(n3450) );
  MUX2IX1 U2420 ( .D0(A[147]), .D1(A[403]), .S(n3181), .Y(n3454) );
  NOR21XL U2421 ( .B(n3455), .A(n3227), .Y(n3449) );
  MUX2IX1 U2422 ( .D0(A[131]), .D1(A[387]), .S(n3181), .Y(n3455) );
  MUX4X1 U2423 ( .D0(n3456), .D1(n3457), .D2(n3458), .D3(n3459), .S0(SH[6]), 
        .S1(SH[5]), .Y(n3431) );
  MUX4X1 U2424 ( .D0(n3460), .D1(n3461), .D2(n3462), .D3(n3463), .S0(n3176), 
        .S1(n3167), .Y(n3459) );
  NOR21XL U2425 ( .B(n3464), .A(n3227), .Y(n3463) );
  MUX2IX1 U2426 ( .D0(A[123]), .D1(A[379]), .S(n3181), .Y(n3464) );
  NOR3XL U2427 ( .A(n3200), .B(n3219), .C(A[363]), .Y(n3462) );
  NOR3XL U2428 ( .A(n3200), .B(n3236), .C(A[371]), .Y(n3461) );
  NOR3XL U2429 ( .A(n3211), .B(n3219), .C(A[355]), .Y(n3460) );
  MUX3X1 U2430 ( .D0(n3465), .D1(n3466), .D2(n3467), .S0(n3170), .S1(n3178), 
        .Y(n3458) );
  NOR4XL U2431 ( .A(n3225), .B(n3188), .C(A[59]), .D(n3172), .Y(n3467) );
  NOR3XL U2432 ( .A(A[43]), .B(n3219), .C(n3190), .Y(n3466) );
  NOR3XL U2433 ( .A(A[35]), .B(n3219), .C(n3190), .Y(n3465) );
  MUX4X1 U2434 ( .D0(n3468), .D1(n3469), .D2(n3470), .D3(n3471), .S0(n3164), 
        .S1(n3177), .Y(n3457) );
  NOR3XL U2435 ( .A(n3202), .B(n3219), .C(A[347]), .Y(n3471) );
  NOR3XL U2436 ( .A(n3202), .B(n3219), .C(A[339]), .Y(n3470) );
  NOR21XL U2437 ( .B(n3472), .A(n3226), .Y(n3469) );
  MUX2IX1 U2438 ( .D0(A[75]), .D1(A[331]), .S(n3181), .Y(n3472) );
  NOR21XL U2439 ( .B(n3473), .A(n3227), .Y(n3468) );
  MUX2IX1 U2440 ( .D0(A[67]), .D1(A[323]), .S(n3180), .Y(n3473) );
  MUX2X1 U2441 ( .D0(n3474), .D1(n3475), .S(n3177), .Y(n3456) );
  NOR4XL U2442 ( .A(n3225), .B(n3188), .C(SH[3]), .D(A[19]), .Y(n3475) );
  MUX2IX1 U2443 ( .D0(n3476), .D1(n3477), .S(n3165), .Y(n3474) );
  NAND2X1 U2444 ( .A(n3478), .B(n3232), .Y(n3477) );
  MUX2IX1 U2445 ( .D0(A[11]), .D1(A[267]), .S(n3180), .Y(n3478) );
  NAND2X1 U2446 ( .A(n3479), .B(n3232), .Y(n3476) );
  MUX2IX1 U2447 ( .D0(A[3]), .D1(A[259]), .S(n3180), .Y(n3479) );
  MUX2IX1 U2448 ( .D0(n3480), .D1(n3481), .S(SH[7]), .Y(B[2]) );
  MUX4X1 U2449 ( .D0(n3482), .D1(n3483), .D2(n3484), .D3(n3485), .S0(SH[5]), 
        .S1(SH[6]), .Y(n3481) );
  MUX4X1 U2450 ( .D0(n3486), .D1(n3487), .D2(n3488), .D3(n3489), .S0(n3176), 
        .S1(n3167), .Y(n3485) );
  NOR3XL U2451 ( .A(A[250]), .B(n3219), .C(n3190), .Y(n3489) );
  NOR3XL U2452 ( .A(A[234]), .B(n3218), .C(n3190), .Y(n3488) );
  NOR3XL U2453 ( .A(A[242]), .B(n3236), .C(n3190), .Y(n3487) );
  NOR3XL U2454 ( .A(A[226]), .B(n3219), .C(n3190), .Y(n3486) );
  MUX4X1 U2455 ( .D0(n3490), .D1(n3491), .D2(n3492), .D3(n3493), .S0(n3176), 
        .S1(n3167), .Y(n3484) );
  NOR3XL U2456 ( .A(A[218]), .B(n3218), .C(n3190), .Y(n3493) );
  AOI21X1 U2457 ( .B(A[202]), .C(n3198), .A(n3214), .Y(n3492) );
  AOI21X1 U2458 ( .B(A[210]), .C(n3198), .A(n3213), .Y(n3491) );
  AOI21X1 U2459 ( .B(A[194]), .C(n3199), .A(n3213), .Y(n3490) );
  MUX4X1 U2460 ( .D0(n3494), .D1(n3495), .D2(n3496), .D3(n3497), .S0(n3174), 
        .S1(n3167), .Y(n3483) );
  NOR3XL U2461 ( .A(A[186]), .B(n3218), .C(n3190), .Y(n3497) );
  NOR3XL U2462 ( .A(A[170]), .B(n3218), .C(n3190), .Y(n3496) );
  NOR3XL U2463 ( .A(A[178]), .B(n3217), .C(n3190), .Y(n3495) );
  NOR3XL U2464 ( .A(A[162]), .B(n3218), .C(n3189), .Y(n3494) );
  MUX4X1 U2465 ( .D0(n3498), .D1(n3499), .D2(n3500), .D3(n3501), .S0(n3176), 
        .S1(n3168), .Y(n3482) );
  NOR3XL U2466 ( .A(A[154]), .B(n3217), .C(n3189), .Y(n3501) );
  NOR21XL U2467 ( .B(n3502), .A(n3229), .Y(n3500) );
  MUX2IX1 U2468 ( .D0(A[138]), .D1(A[394]), .S(n3183), .Y(n3502) );
  NOR21XL U2469 ( .B(n3503), .A(n3228), .Y(n3499) );
  MUX2IX1 U2470 ( .D0(A[146]), .D1(A[402]), .S(n3180), .Y(n3503) );
  NOR21XL U2471 ( .B(n3504), .A(n3228), .Y(n3498) );
  MUX2IX1 U2472 ( .D0(A[130]), .D1(A[386]), .S(n3180), .Y(n3504) );
  MUX4X1 U2473 ( .D0(n3505), .D1(n3506), .D2(n3507), .D3(n3508), .S0(SH[6]), 
        .S1(n3163), .Y(n3480) );
  MUX4X1 U2474 ( .D0(n3509), .D1(n3510), .D2(n3511), .D3(n3512), .S0(n3176), 
        .S1(n3167), .Y(n3508) );
  NOR21XL U2475 ( .B(n3513), .A(n3227), .Y(n3512) );
  MUX2IX1 U2476 ( .D0(A[122]), .D1(A[378]), .S(n3180), .Y(n3513) );
  NOR3XL U2477 ( .A(n3201), .B(n3217), .C(A[362]), .Y(n3511) );
  NOR3XL U2478 ( .A(n3203), .B(n3218), .C(A[370]), .Y(n3510) );
  NOR3XL U2479 ( .A(n3204), .B(n3217), .C(A[354]), .Y(n3509) );
  MUX3X1 U2480 ( .D0(n3514), .D1(n3515), .D2(n3516), .S0(n3169), .S1(SH[4]), 
        .Y(n3507) );
  NOR4XL U2481 ( .A(n3225), .B(n3188), .C(A[58]), .D(n3172), .Y(n3516) );
  NOR3XL U2482 ( .A(A[42]), .B(n3217), .C(n3189), .Y(n3515) );
  NOR3XL U2483 ( .A(A[34]), .B(n3218), .C(n3189), .Y(n3514) );
  MUX4X1 U2484 ( .D0(n3517), .D1(n3518), .D2(n3519), .D3(n3520), .S0(n3164), 
        .S1(n3177), .Y(n3506) );
  NOR3XL U2485 ( .A(n3211), .B(n3216), .C(A[346]), .Y(n3520) );
  NOR3XL U2486 ( .A(n3211), .B(n3216), .C(A[338]), .Y(n3519) );
  NOR21XL U2487 ( .B(n3521), .A(n3227), .Y(n3518) );
  MUX2IX1 U2488 ( .D0(A[74]), .D1(A[330]), .S(n3180), .Y(n3521) );
  NOR21XL U2489 ( .B(n3522), .A(n3228), .Y(n3517) );
  MUX2IX1 U2490 ( .D0(A[66]), .D1(A[322]), .S(n3180), .Y(n3522) );
  MUX2X1 U2491 ( .D0(n3523), .D1(n3524), .S(n3177), .Y(n3505) );
  NOR4XL U2492 ( .A(n3225), .B(n3188), .C(n3170), .D(A[18]), .Y(n3524) );
  MUX2IX1 U2493 ( .D0(n3525), .D1(n3526), .S(n3164), .Y(n3523) );
  NAND2X1 U2494 ( .A(n3527), .B(n3234), .Y(n3526) );
  MUX2IX1 U2495 ( .D0(A[10]), .D1(A[266]), .S(n3180), .Y(n3527) );
  NAND2X1 U2496 ( .A(n3528), .B(n3233), .Y(n3525) );
  MUX2IX1 U2497 ( .D0(A[2]), .D1(A[258]), .S(n3181), .Y(n3528) );
  MUX2IX1 U2498 ( .D0(n3529), .D1(n3530), .S(SH[7]), .Y(B[1]) );
  MUX4X1 U2499 ( .D0(n3531), .D1(n3532), .D2(n3533), .D3(n3534), .S0(SH[5]), 
        .S1(n3162), .Y(n3530) );
  MUX4X1 U2500 ( .D0(n3535), .D1(n3536), .D2(n3537), .D3(n3538), .S0(n3176), 
        .S1(n3168), .Y(n3534) );
  NOR3XL U2501 ( .A(A[249]), .B(n3217), .C(n3193), .Y(n3538) );
  NOR3XL U2502 ( .A(A[233]), .B(n3220), .C(n3209), .Y(n3537) );
  NOR3XL U2503 ( .A(A[241]), .B(n3216), .C(n3189), .Y(n3536) );
  NOR3XL U2504 ( .A(A[225]), .B(n3218), .C(SH[8]), .Y(n3535) );
  MUX4X1 U2505 ( .D0(n3539), .D1(n3540), .D2(n3541), .D3(n3542), .S0(n3176), 
        .S1(n3168), .Y(n3533) );
  NOR3XL U2506 ( .A(A[217]), .B(n3218), .C(n3193), .Y(n3542) );
  NOR21XL U2507 ( .B(n3543), .A(n3228), .Y(n3541) );
  MUX2IX1 U2508 ( .D0(A[201]), .D1(A[457]), .S(n3181), .Y(n3543) );
  NOR21XL U2509 ( .B(n3544), .A(n3229), .Y(n3540) );
  MUX2IX1 U2510 ( .D0(A[209]), .D1(A[465]), .S(n3181), .Y(n3544) );
  NOR21XL U2511 ( .B(n3545), .A(n3229), .Y(n3539) );
  MUX2IX1 U2512 ( .D0(A[193]), .D1(A[449]), .S(n3181), .Y(n3545) );
  MUX4X1 U2513 ( .D0(n3546), .D1(n3547), .D2(n3548), .D3(n3549), .S0(n3175), 
        .S1(n3167), .Y(n3532) );
  NOR3XL U2514 ( .A(A[185]), .B(n3216), .C(n3189), .Y(n3549) );
  NOR3XL U2515 ( .A(A[169]), .B(n3216), .C(n3209), .Y(n3548) );
  NOR3XL U2516 ( .A(A[177]), .B(n3215), .C(n3207), .Y(n3547) );
  NOR3XL U2517 ( .A(A[161]), .B(n3217), .C(n3207), .Y(n3546) );
  MUX4X1 U2518 ( .D0(n3550), .D1(n3551), .D2(n3552), .D3(n3553), .S0(n3175), 
        .S1(n3168), .Y(n3531) );
  NOR3XL U2519 ( .A(A[153]), .B(n3215), .C(n3209), .Y(n3553) );
  NOR21XL U2520 ( .B(n3554), .A(n3230), .Y(n3552) );
  MUX2IX1 U2521 ( .D0(A[137]), .D1(A[393]), .S(n3182), .Y(n3554) );
  NOR21XL U2522 ( .B(n3555), .A(n3228), .Y(n3551) );
  MUX2IX1 U2523 ( .D0(A[145]), .D1(A[401]), .S(n3182), .Y(n3555) );
  NOR21XL U2524 ( .B(n3556), .A(n3228), .Y(n3550) );
  MUX2IX1 U2525 ( .D0(A[129]), .D1(A[385]), .S(n3182), .Y(n3556) );
  MUX4X1 U2526 ( .D0(n3557), .D1(n3558), .D2(n3559), .D3(n3560), .S0(SH[6]), 
        .S1(n3163), .Y(n3529) );
  MUX4X1 U2527 ( .D0(n3561), .D1(n3562), .D2(n3563), .D3(n3564), .S0(n3175), 
        .S1(n3169), .Y(n3560) );
  NOR21XL U2528 ( .B(n3565), .A(n3229), .Y(n3564) );
  MUX2IX1 U2529 ( .D0(A[121]), .D1(A[377]), .S(n3183), .Y(n3565) );
  NOR3XL U2530 ( .A(n3212), .B(n3215), .C(A[361]), .Y(n3563) );
  NOR3XL U2531 ( .A(n3203), .B(n3217), .C(A[369]), .Y(n3562) );
  NOR3XL U2532 ( .A(n3201), .B(n3215), .C(A[353]), .Y(n3561) );
  MUX3X1 U2533 ( .D0(n3566), .D1(n3567), .D2(n3568), .S0(n3170), .S1(n3178), 
        .Y(n3559) );
  NOR4XL U2534 ( .A(n3225), .B(n3187), .C(A[57]), .D(n3172), .Y(n3568) );
  NOR3XL U2535 ( .A(A[41]), .B(n3215), .C(n3209), .Y(n3567) );
  NOR3XL U2536 ( .A(A[33]), .B(n3218), .C(SH[8]), .Y(n3566) );
  MUX4X1 U2537 ( .D0(n3569), .D1(n3570), .D2(n3571), .D3(n3572), .S0(n3164), 
        .S1(n3176), .Y(n3558) );
  NOR3XL U2538 ( .A(n3201), .B(n3215), .C(A[345]), .Y(n3572) );
  NOR3XL U2539 ( .A(n3200), .B(n3215), .C(A[337]), .Y(n3571) );
  NOR21XL U2540 ( .B(n3573), .A(n3230), .Y(n3570) );
  MUX2IX1 U2541 ( .D0(A[73]), .D1(A[329]), .S(n3183), .Y(n3573) );
  NOR21XL U2542 ( .B(n3574), .A(n3229), .Y(n3569) );
  MUX2IX1 U2543 ( .D0(A[65]), .D1(A[321]), .S(n3183), .Y(n3574) );
  MUX2X1 U2544 ( .D0(n3575), .D1(n3576), .S(n3177), .Y(n3557) );
  NOR4XL U2545 ( .A(n3226), .B(n3188), .C(n3170), .D(A[17]), .Y(n3576) );
  MUX2IX1 U2546 ( .D0(n3577), .D1(n3578), .S(n3164), .Y(n3575) );
  NAND2X1 U2547 ( .A(n3579), .B(n3234), .Y(n3578) );
  MUX2IX1 U2548 ( .D0(A[9]), .D1(A[265]), .S(n3183), .Y(n3579) );
  NAND2X1 U2549 ( .A(n3580), .B(n3233), .Y(n3577) );
  MUX2IX1 U2550 ( .D0(A[1]), .D1(A[257]), .S(n3183), .Y(n3580) );
  MUX2IX1 U2551 ( .D0(n3581), .D1(n3582), .S(SH[7]), .Y(B[0]) );
  MUX4X1 U2552 ( .D0(n3583), .D1(n3584), .D2(n3585), .D3(n3586), .S0(SH[5]), 
        .S1(n3162), .Y(n3582) );
  MUX4X1 U2553 ( .D0(n3587), .D1(n3588), .D2(n3589), .D3(n3590), .S0(n3174), 
        .S1(n3168), .Y(n3586) );
  NOR3XL U2554 ( .A(A[248]), .B(n3216), .C(SH[8]), .Y(n3590) );
  NOR3XL U2555 ( .A(A[232]), .B(n3217), .C(n3209), .Y(n3589) );
  NOR3XL U2556 ( .A(A[240]), .B(n3237), .C(SH[8]), .Y(n3588) );
  NOR3XL U2557 ( .A(A[224]), .B(n3216), .C(n3209), .Y(n3587) );
  MUX4X1 U2558 ( .D0(n3591), .D1(n3592), .D2(n3593), .D3(n3594), .S0(n3174), 
        .S1(n3169), .Y(n3585) );
  NOR3XL U2559 ( .A(A[216]), .B(SH[9]), .C(n3208), .Y(n3594) );
  NOR21XL U2560 ( .B(n3595), .A(n3229), .Y(n3593) );
  MUX2IX1 U2561 ( .D0(A[200]), .D1(A[456]), .S(n3184), .Y(n3595) );
  NOR21XL U2562 ( .B(n3596), .A(n3230), .Y(n3592) );
  MUX2IX1 U2563 ( .D0(A[208]), .D1(A[464]), .S(n3184), .Y(n3596) );
  NOR21XL U2564 ( .B(n3597), .A(n3230), .Y(n3591) );
  MUX2IX1 U2565 ( .D0(A[192]), .D1(A[448]), .S(n3184), .Y(n3597) );
  MUX4X1 U2566 ( .D0(n3598), .D1(n3599), .D2(n3600), .D3(n3601), .S0(n3173), 
        .S1(n3168), .Y(n3584) );
  NOR3XL U2567 ( .A(A[184]), .B(n3216), .C(n3209), .Y(n3601) );
  NOR3XL U2568 ( .A(A[168]), .B(n3216), .C(SH[8]), .Y(n3600) );
  NOR3XL U2569 ( .A(A[176]), .B(n3236), .C(SH[8]), .Y(n3599) );
  NOR3XL U2570 ( .A(A[160]), .B(n3236), .C(n3189), .Y(n3598) );
  MUX4X1 U2571 ( .D0(n3602), .D1(n3603), .D2(n3604), .D3(n3605), .S0(n3173), 
        .S1(n3168), .Y(n3583) );
  NOR3XL U2572 ( .A(A[152]), .B(n3216), .C(SH[8]), .Y(n3605) );
  NOR21XL U2573 ( .B(n3606), .A(n3231), .Y(n3604) );
  MUX2IX1 U2574 ( .D0(A[136]), .D1(A[392]), .S(n3186), .Y(n3606) );
  NOR21XL U2575 ( .B(n3607), .A(n3230), .Y(n3603) );
  MUX2IX1 U2576 ( .D0(A[144]), .D1(A[400]), .S(n3185), .Y(n3607) );
  NOR21XL U2577 ( .B(n3608), .A(n3231), .Y(n3602) );
  MUX2IX1 U2578 ( .D0(A[128]), .D1(A[384]), .S(n3185), .Y(n3608) );
  MUX4X1 U2579 ( .D0(n3609), .D1(n3610), .D2(n3611), .D3(n3612), .S0(SH[6]), 
        .S1(n3163), .Y(n3581) );
  MUX4X1 U2580 ( .D0(n3613), .D1(n3614), .D2(n3615), .D3(n3616), .S0(n3173), 
        .S1(n3168), .Y(n3612) );
  NOR21XL U2581 ( .B(n3617), .A(n3231), .Y(n3616) );
  MUX2IX1 U2582 ( .D0(A[120]), .D1(A[376]), .S(n3186), .Y(n3617) );
  NOR3XL U2583 ( .A(n3201), .B(SH[9]), .C(A[360]), .Y(n3615) );
  NOR3XL U2584 ( .A(n3202), .B(n3217), .C(A[368]), .Y(n3614) );
  NOR3XL U2585 ( .A(n3202), .B(n3215), .C(A[352]), .Y(n3613) );
  MUX3X1 U2586 ( .D0(n3618), .D1(n3619), .D2(n3620), .S0(n3170), .S1(SH[4]), 
        .Y(n3611) );
  NOR4XL U2587 ( .A(n3226), .B(n3188), .C(A[56]), .D(n3172), .Y(n3620) );
  NOR3XL U2588 ( .A(A[40]), .B(SH[9]), .C(n3209), .Y(n3619) );
  NOR3XL U2589 ( .A(A[32]), .B(n3215), .C(n3189), .Y(n3618) );
  MUX4X1 U2590 ( .D0(n3621), .D1(n3622), .D2(n3623), .D3(n3624), .S0(n3164), 
        .S1(n3176), .Y(n3610) );
  NOR3XL U2591 ( .A(n3199), .B(n3236), .C(A[344]), .Y(n3624) );
  NOR3XL U2592 ( .A(n3211), .B(SH[9]), .C(A[336]), .Y(n3623) );
  NOR21XL U2593 ( .B(n3625), .A(n3231), .Y(n3622) );
  MUX2IX1 U2594 ( .D0(A[72]), .D1(A[328]), .S(n3186), .Y(n3625) );
  NOR21XL U2595 ( .B(n3626), .A(n3231), .Y(n3621) );
  MUX2IX1 U2596 ( .D0(A[64]), .D1(A[320]), .S(n3186), .Y(n3626) );
  MUX2X1 U2597 ( .D0(n3627), .D1(n3628), .S(n3177), .Y(n3609) );
  NOR4XL U2598 ( .A(n3225), .B(n3188), .C(SH[3]), .D(A[16]), .Y(n3628) );
  MUX2IX1 U2599 ( .D0(n3629), .D1(n3630), .S(n3165), .Y(n3627) );
  NAND2X1 U2600 ( .A(n3631), .B(n3232), .Y(n3630) );
  MUX2IX1 U2601 ( .D0(A[8]), .D1(A[264]), .S(n3186), .Y(n3631) );
  NAND2X1 U2602 ( .A(n3632), .B(n3233), .Y(n3629) );
  MUX2IX1 U2603 ( .D0(A[0]), .D1(A[256]), .S(n3180), .Y(n3632) );
endmodule


module SNPS_CLOCK_GATE_HIGH_regx_a0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module dbnc_a0_0 ( o_dbc, o_chg, i_org, clk, rstz );
  input i_org, clk, rstz;
  output o_dbc, o_chg;
  wire   d_org_0_, N16, N17, N18, N19, N20, net8993, n5, n6, n7, n8, n9, n10,
         n11, n12, n1, n2, n3, n4;
  wire   [3:0] db_cnt;

  SNPS_CLOCK_GATE_HIGH_dbnc_a0_0 clk_gate_db_cnt_reg ( .CLK(clk), .EN(N16), 
        .ENCLK(net8993), .TE(1'b0) );
  DFFRQX1 d_org_reg_0_ ( .D(i_org), .C(clk), .XR(rstz), .Q(d_org_0_) );
  DFFRQX1 db_cnt_reg_3_ ( .D(N20), .C(net8993), .XR(rstz), .Q(db_cnt[3]) );
  DFFRQX1 db_cnt_reg_2_ ( .D(N19), .C(net8993), .XR(rstz), .Q(db_cnt[2]) );
  DFFRQX1 db_cnt_reg_1_ ( .D(N18), .C(net8993), .XR(rstz), .Q(db_cnt[1]) );
  DFFRQX1 db_cnt_reg_0_ ( .D(N17), .C(net8993), .XR(rstz), .Q(db_cnt[0]) );
  DFFRQX1 d_org_reg_1_ ( .D(n12), .C(net8993), .XR(rstz), .Q(o_dbc) );
  INVX1 U3 ( .A(n8), .Y(n1) );
  NOR2X1 U4 ( .A(n6), .B(n5), .Y(n8) );
  NOR2X1 U5 ( .A(n3), .B(n7), .Y(n5) );
  OAI22X1 U6 ( .A(n1), .B(n3), .C(n7), .D(n1), .Y(N20) );
  NOR2X1 U7 ( .A(n10), .B(n1), .Y(N18) );
  XNOR2XL U8 ( .A(n4), .B(n2), .Y(n10) );
  GEN2XL U9 ( .D(n8), .E(n4), .C(N17), .B(db_cnt[2]), .A(n9), .Y(N19) );
  NOR4XL U10 ( .A(db_cnt[2]), .B(n2), .C(n4), .D(n1), .Y(n9) );
  NAND3X1 U11 ( .A(db_cnt[1]), .B(db_cnt[0]), .C(db_cnt[2]), .Y(n7) );
  NOR2X1 U12 ( .A(n1), .B(db_cnt[0]), .Y(N17) );
  XNOR2XL U13 ( .A(o_dbc), .B(d_org_0_), .Y(n6) );
  AO22AXL U14 ( .A(d_org_0_), .B(o_chg), .C(o_dbc), .D(o_chg), .Y(n12) );
  NOR21XL U15 ( .B(n5), .A(n6), .Y(o_chg) );
  INVX1 U16 ( .A(db_cnt[3]), .Y(n3) );
  INVX1 U17 ( .A(db_cnt[0]), .Y(n2) );
  INVX1 U18 ( .A(db_cnt[1]), .Y(n4) );
  NAND3X1 U19 ( .A(n6), .B(n2), .C(n11), .Y(N16) );
  NOR3XL U20 ( .A(db_cnt[1]), .B(db_cnt[3]), .C(db_cnt[2]), .Y(n11) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dbnc_a0_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module dbnc_a0_1 ( o_dbc, o_chg, i_org, clk, rstz );
  input i_org, clk, rstz;
  output o_dbc, o_chg;
  wire   d_org_0_, N16, N17, N18, N19, N20, net9011, n5, n6, n7, n8, n9, n10,
         n11, n12, n1, n2, n3, n4;
  wire   [3:0] db_cnt;

  SNPS_CLOCK_GATE_HIGH_dbnc_a0_1 clk_gate_db_cnt_reg ( .CLK(clk), .EN(N16), 
        .ENCLK(net9011), .TE(1'b0) );
  DFFRQX1 d_org_reg_0_ ( .D(i_org), .C(clk), .XR(rstz), .Q(d_org_0_) );
  DFFRQX1 db_cnt_reg_3_ ( .D(N20), .C(net9011), .XR(rstz), .Q(db_cnt[3]) );
  DFFRQX1 db_cnt_reg_2_ ( .D(N19), .C(net9011), .XR(rstz), .Q(db_cnt[2]) );
  DFFRQX1 db_cnt_reg_1_ ( .D(N18), .C(net9011), .XR(rstz), .Q(db_cnt[1]) );
  DFFRQX1 db_cnt_reg_0_ ( .D(N17), .C(net9011), .XR(rstz), .Q(db_cnt[0]) );
  DFFRQX1 d_org_reg_1_ ( .D(n12), .C(net9011), .XR(rstz), .Q(o_dbc) );
  INVX1 U3 ( .A(n8), .Y(n1) );
  NOR2X1 U4 ( .A(n6), .B(n5), .Y(n8) );
  NOR2X1 U5 ( .A(n3), .B(n7), .Y(n5) );
  OAI22X1 U6 ( .A(n1), .B(n3), .C(n7), .D(n1), .Y(N20) );
  NOR2X1 U7 ( .A(n10), .B(n1), .Y(N18) );
  XNOR2XL U8 ( .A(n4), .B(n2), .Y(n10) );
  GEN2XL U9 ( .D(n8), .E(n4), .C(N17), .B(db_cnt[2]), .A(n9), .Y(N19) );
  NOR4XL U10 ( .A(db_cnt[2]), .B(n2), .C(n4), .D(n1), .Y(n9) );
  NAND3X1 U11 ( .A(db_cnt[1]), .B(db_cnt[0]), .C(db_cnt[2]), .Y(n7) );
  NOR2X1 U12 ( .A(n1), .B(db_cnt[0]), .Y(N17) );
  XNOR2XL U13 ( .A(o_dbc), .B(d_org_0_), .Y(n6) );
  AO22AXL U14 ( .A(d_org_0_), .B(o_chg), .C(o_dbc), .D(o_chg), .Y(n12) );
  NOR21XL U15 ( .B(n5), .A(n6), .Y(o_chg) );
  INVX1 U16 ( .A(db_cnt[3]), .Y(n3) );
  INVX1 U17 ( .A(db_cnt[0]), .Y(n2) );
  INVX1 U18 ( .A(db_cnt[1]), .Y(n4) );
  NAND3X1 U19 ( .A(n6), .B(n2), .C(n11), .Y(N16) );
  NOR3XL U20 ( .A(db_cnt[1]), .B(db_cnt[3]), .C(db_cnt[2]), .Y(n11) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dbnc_a0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module dbnc_WIDTH2_TIMEOUT2_0 ( o_dbc, o_chg, i_org, clk, rstz );
  input i_org, clk, rstz;
  output o_dbc, o_chg;
  wire   d_org_0_, n1, n7, n8, n9, n10, n11;
  wire   [1:0] db_cnt;

  DFFRQX1 db_cnt_reg_1_ ( .D(n8), .C(clk), .XR(rstz), .Q(db_cnt[1]) );
  DFFRQX1 db_cnt_reg_0_ ( .D(n7), .C(clk), .XR(rstz), .Q(db_cnt[0]) );
  DFFRQX1 d_org_reg_0_ ( .D(i_org), .C(clk), .XR(rstz), .Q(d_org_0_) );
  DFFRQX1 d_org_reg_1_ ( .D(n9), .C(clk), .XR(rstz), .Q(o_dbc) );
  XNOR2XL U3 ( .A(n1), .B(d_org_0_), .Y(n11) );
  ENOX1 U4 ( .A(o_chg), .B(n1), .C(d_org_0_), .D(o_chg), .Y(n9) );
  NOR32XL U5 ( .B(n11), .C(db_cnt[1]), .A(db_cnt[0]), .Y(o_chg) );
  INVX1 U6 ( .A(o_dbc), .Y(n1) );
  NAND21X1 U7 ( .B(db_cnt[1]), .A(n11), .Y(n10) );
  NOR21XL U8 ( .B(db_cnt[0]), .A(n10), .Y(n8) );
  NOR2X1 U9 ( .A(db_cnt[0]), .B(n10), .Y(n7) );
endmodule


module dbnc_WIDTH2_TIMEOUT2_1 ( o_dbc, o_chg, i_org, clk, rstz );
  input i_org, clk, rstz;
  output o_dbc, o_chg;
  wire   d_org_0_, n1, n7, n8, n9, n10, n11;
  wire   [1:0] db_cnt;

  DFFRQX1 db_cnt_reg_1_ ( .D(n8), .C(clk), .XR(rstz), .Q(db_cnt[1]) );
  DFFRQX1 db_cnt_reg_0_ ( .D(n7), .C(clk), .XR(rstz), .Q(db_cnt[0]) );
  DFFRQX1 d_org_reg_0_ ( .D(i_org), .C(clk), .XR(rstz), .Q(d_org_0_) );
  DFFRQX1 d_org_reg_1_ ( .D(n9), .C(clk), .XR(rstz), .Q(o_dbc) );
  XNOR2XL U3 ( .A(n1), .B(d_org_0_), .Y(n11) );
  ENOX1 U4 ( .A(o_chg), .B(n1), .C(d_org_0_), .D(o_chg), .Y(n9) );
  NOR32XL U5 ( .B(n11), .C(db_cnt[1]), .A(db_cnt[0]), .Y(o_chg) );
  INVX1 U6 ( .A(o_dbc), .Y(n1) );
  NAND21X1 U7 ( .B(db_cnt[1]), .A(n11), .Y(n10) );
  NOR21XL U8 ( .B(db_cnt[0]), .A(n10), .Y(n8) );
  NOR2X1 U9 ( .A(db_cnt[0]), .B(n10), .Y(n7) );
endmodule


module dbnc_WIDTH2_TIMEOUT2_2 ( o_dbc, o_chg, i_org, clk, rstz );
  input i_org, clk, rstz;
  output o_dbc, o_chg;
  wire   d_org_0_, n1, n7, n8, n9, n10, n11;
  wire   [1:0] db_cnt;

  DFFRQX1 db_cnt_reg_1_ ( .D(n8), .C(clk), .XR(rstz), .Q(db_cnt[1]) );
  DFFRQX1 db_cnt_reg_0_ ( .D(n7), .C(clk), .XR(rstz), .Q(db_cnt[0]) );
  DFFRQX1 d_org_reg_0_ ( .D(i_org), .C(clk), .XR(rstz), .Q(d_org_0_) );
  DFFRQX1 d_org_reg_1_ ( .D(n9), .C(clk), .XR(rstz), .Q(o_dbc) );
  XNOR2XL U3 ( .A(n1), .B(d_org_0_), .Y(n11) );
  ENOX1 U4 ( .A(o_chg), .B(n1), .C(d_org_0_), .D(o_chg), .Y(n9) );
  NOR32XL U5 ( .B(n11), .C(db_cnt[1]), .A(db_cnt[0]), .Y(o_chg) );
  INVX1 U6 ( .A(o_dbc), .Y(n1) );
  NAND21X1 U7 ( .B(db_cnt[1]), .A(n11), .Y(n10) );
  NOR21XL U8 ( .B(db_cnt[0]), .A(n10), .Y(n8) );
  NOR2X1 U9 ( .A(db_cnt[0]), .B(n10), .Y(n7) );
endmodule


module dbnc_WIDTH2_TIMEOUT2_3 ( o_dbc, o_chg, i_org, clk, rstz );
  input i_org, clk, rstz;
  output o_dbc, o_chg;
  wire   d_org_0_, n1, n7, n8, n9, n10, n11;
  wire   [1:0] db_cnt;

  DFFRQX1 db_cnt_reg_1_ ( .D(n8), .C(clk), .XR(rstz), .Q(db_cnt[1]) );
  DFFRQX1 db_cnt_reg_0_ ( .D(n7), .C(clk), .XR(rstz), .Q(db_cnt[0]) );
  DFFRQX1 d_org_reg_0_ ( .D(i_org), .C(clk), .XR(rstz), .Q(d_org_0_) );
  DFFRQX1 d_org_reg_1_ ( .D(n9), .C(clk), .XR(rstz), .Q(o_dbc) );
  XNOR2XL U3 ( .A(n1), .B(d_org_0_), .Y(n11) );
  ENOX1 U4 ( .A(o_chg), .B(n1), .C(d_org_0_), .D(o_chg), .Y(n9) );
  NOR32XL U5 ( .B(n11), .C(db_cnt[1]), .A(db_cnt[0]), .Y(o_chg) );
  INVX1 U6 ( .A(o_dbc), .Y(n1) );
  NAND21X1 U7 ( .B(db_cnt[1]), .A(n11), .Y(n10) );
  NOR21XL U8 ( .B(db_cnt[0]), .A(n10), .Y(n8) );
  NOR2X1 U9 ( .A(db_cnt[0]), .B(n10), .Y(n7) );
endmodule


module dbnc_WIDTH2_TIMEOUT2_4 ( o_dbc, o_chg, i_org, clk, rstz );
  input i_org, clk, rstz;
  output o_dbc, o_chg;
  wire   d_org_0_, n1, n7, n8, n9, n10, n11;
  wire   [1:0] db_cnt;

  DFFRQX1 db_cnt_reg_1_ ( .D(n8), .C(clk), .XR(rstz), .Q(db_cnt[1]) );
  DFFRQX1 db_cnt_reg_0_ ( .D(n7), .C(clk), .XR(rstz), .Q(db_cnt[0]) );
  DFFRQX1 d_org_reg_0_ ( .D(i_org), .C(clk), .XR(rstz), .Q(d_org_0_) );
  DFFRQX1 d_org_reg_1_ ( .D(n9), .C(clk), .XR(rstz), .Q(o_dbc) );
  XNOR2XL U3 ( .A(n1), .B(d_org_0_), .Y(n11) );
  ENOX1 U4 ( .A(o_chg), .B(n1), .C(d_org_0_), .D(o_chg), .Y(n9) );
  NOR32XL U5 ( .B(n11), .C(db_cnt[1]), .A(db_cnt[0]), .Y(o_chg) );
  INVX1 U6 ( .A(o_dbc), .Y(n1) );
  NAND21X1 U7 ( .B(db_cnt[1]), .A(n11), .Y(n10) );
  NOR21XL U8 ( .B(db_cnt[0]), .A(n10), .Y(n8) );
  NOR2X1 U9 ( .A(db_cnt[0]), .B(n10), .Y(n7) );
endmodule


module dbnc_WIDTH2_TIMEOUT2_5 ( o_dbc, o_chg, i_org, clk, rstz );
  input i_org, clk, rstz;
  output o_dbc, o_chg;
  wire   d_org_0_, n1, n7, n8, n9, n10, n11;
  wire   [1:0] db_cnt;

  DFFRQX1 db_cnt_reg_1_ ( .D(n8), .C(clk), .XR(rstz), .Q(db_cnt[1]) );
  DFFRQX1 db_cnt_reg_0_ ( .D(n7), .C(clk), .XR(rstz), .Q(db_cnt[0]) );
  DFFRQX1 d_org_reg_0_ ( .D(i_org), .C(clk), .XR(rstz), .Q(d_org_0_) );
  DFFRQX1 d_org_reg_1_ ( .D(n9), .C(clk), .XR(rstz), .Q(o_dbc) );
  XNOR2XL U3 ( .A(n1), .B(d_org_0_), .Y(n11) );
  ENOX1 U4 ( .A(o_chg), .B(n1), .C(d_org_0_), .D(o_chg), .Y(n9) );
  NOR32XL U5 ( .B(n11), .C(db_cnt[1]), .A(db_cnt[0]), .Y(o_chg) );
  INVX1 U6 ( .A(o_dbc), .Y(n1) );
  NAND21X1 U7 ( .B(db_cnt[1]), .A(n11), .Y(n10) );
  NOR21XL U8 ( .B(db_cnt[0]), .A(n10), .Y(n8) );
  NOR2X1 U9 ( .A(db_cnt[0]), .B(n10), .Y(n7) );
endmodule


module dbnc_WIDTH2_TIMEOUT2_6 ( o_dbc, o_chg, i_org, clk, rstz );
  input i_org, clk, rstz;
  output o_dbc, o_chg;
  wire   d_org_0_, n1, n7, n8, n9, n10, n11;
  wire   [1:0] db_cnt;

  DFFRQX1 db_cnt_reg_1_ ( .D(n8), .C(clk), .XR(rstz), .Q(db_cnt[1]) );
  DFFRQX1 db_cnt_reg_0_ ( .D(n7), .C(clk), .XR(rstz), .Q(db_cnt[0]) );
  DFFRQX1 d_org_reg_0_ ( .D(i_org), .C(clk), .XR(rstz), .Q(d_org_0_) );
  DFFRQX1 d_org_reg_1_ ( .D(n9), .C(clk), .XR(rstz), .Q(o_dbc) );
  XNOR2XL U3 ( .A(n1), .B(d_org_0_), .Y(n11) );
  ENOX1 U4 ( .A(o_chg), .B(n1), .C(d_org_0_), .D(o_chg), .Y(n9) );
  NOR32XL U5 ( .B(n11), .C(db_cnt[1]), .A(db_cnt[0]), .Y(o_chg) );
  INVX1 U6 ( .A(o_dbc), .Y(n1) );
  NAND21X1 U7 ( .B(db_cnt[1]), .A(n11), .Y(n10) );
  NOR21XL U8 ( .B(db_cnt[0]), .A(n10), .Y(n8) );
  NOR2X1 U9 ( .A(db_cnt[0]), .B(n10), .Y(n7) );
endmodule


module glreg_a0_7 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net9029;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_7 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9029), .TE(1'b0) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net9029), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net9029), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net9029), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net9029), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net9029), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net9029), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net9029), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net9029), .XR(arstz), .Q(rdat[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_7 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_8 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net9047;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_8 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9047), .TE(1'b0) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net9047), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net9047), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net9047), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net9047), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net9047), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net9047), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net9047), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net9047), .XR(arstz), .Q(rdat[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_8 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_9 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net9065;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_9 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9065), .TE(1'b0) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net9065), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net9065), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net9065), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net9065), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net9065), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net9065), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net9065), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net9065), .XR(arstz), .Q(rdat[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_9 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_WIDTH1_1 ( clk, arstz, we, wdat, rdat );
  input [0:0] wdat;
  output [0:0] rdat;
  input clk, arstz, we;
  wire   n2;

  DFFRQX1 mem_reg_0_ ( .D(n2), .C(clk), .XR(arstz), .Q(rdat[0]) );
  AO22AXL U2 ( .A(we), .B(wdat[0]), .C(rdat[0]), .D(we), .Y(n2) );
endmodule


module glreg_WIDTH7_0 ( clk, arstz, we, wdat, rdat );
  input [6:0] wdat;
  output [6:0] rdat;
  input clk, arstz, we;
  wire   net9083;

  SNPS_CLOCK_GATE_HIGH_glreg_WIDTH7_0 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9083), .TE(1'b0) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net9083), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net9083), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net9083), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net9083), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net9083), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net9083), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net9083), .XR(arstz), .Q(rdat[6]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_WIDTH7_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module dbnc_WIDTH2_TIMEOUT2_7 ( o_dbc, o_chg, i_org, clk, rstz );
  input i_org, clk, rstz;
  output o_dbc, o_chg;
  wire   d_org_0_, n1, n7, n8, n9, n10, n11;
  wire   [1:0] db_cnt;

  DFFRQX1 db_cnt_reg_1_ ( .D(n8), .C(clk), .XR(rstz), .Q(db_cnt[1]) );
  DFFRQX1 db_cnt_reg_0_ ( .D(n7), .C(clk), .XR(rstz), .Q(db_cnt[0]) );
  DFFRQX1 d_org_reg_0_ ( .D(i_org), .C(clk), .XR(rstz), .Q(d_org_0_) );
  DFFRQX1 d_org_reg_1_ ( .D(n9), .C(clk), .XR(rstz), .Q(o_dbc) );
  XNOR2XL U3 ( .A(n1), .B(d_org_0_), .Y(n11) );
  ENOX1 U4 ( .A(o_chg), .B(n1), .C(d_org_0_), .D(o_chg), .Y(n9) );
  NOR32XL U5 ( .B(n11), .C(db_cnt[1]), .A(db_cnt[0]), .Y(o_chg) );
  INVX1 U6 ( .A(o_dbc), .Y(n1) );
  NAND21X1 U7 ( .B(db_cnt[1]), .A(n11), .Y(n10) );
  NOR21XL U8 ( .B(db_cnt[0]), .A(n10), .Y(n8) );
  NOR2X1 U9 ( .A(db_cnt[0]), .B(n10), .Y(n7) );
endmodule


module glreg_a0_10 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net9101;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_10 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9101), .TE(1'b0) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net9101), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net9101), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net9101), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net9101), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net9101), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net9101), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net9101), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net9101), .XR(arstz), .Q(rdat[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_10 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_11 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net9119;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_11 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9119), .TE(1'b0) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net9119), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net9119), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net9119), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net9119), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net9119), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net9119), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net9119), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net9119), .XR(arstz), .Q(rdat[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_11 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_12 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net9137;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_12 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9137), .TE(1'b0) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net9137), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net9137), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net9137), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net9137), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net9137), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net9137), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net9137), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net9137), .XR(arstz), .Q(rdat[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_12 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_13 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net9155;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_13 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9155), .TE(1'b0) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net9155), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net9155), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net9155), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net9155), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net9155), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net9155), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net9155), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net9155), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_13 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_14 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net9173;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_14 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9173), .TE(1'b0) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net9173), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net9173), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net9173), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net9173), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net9173), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net9173), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net9173), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net9173), .XR(arstz), .Q(rdat[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_14 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_WIDTH6_0 ( clk, arstz, we, wdat, rdat );
  input [5:0] wdat;
  output [5:0] rdat;
  input clk, arstz, we;
  wire   net9191;

  SNPS_CLOCK_GATE_HIGH_glreg_WIDTH6_0 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9191), .TE(1'b0) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net9191), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net9191), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net9191), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net9191), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net9191), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net9191), .XR(arstz), .Q(rdat[2]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_WIDTH6_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_WIDTH6_1 ( clk, arstz, we, wdat, rdat );
  input [5:0] wdat;
  output [5:0] rdat;
  input clk, arstz, we;
  wire   net9209;

  SNPS_CLOCK_GATE_HIGH_glreg_WIDTH6_1 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9209), .TE(1'b0) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net9209), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net9209), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net9209), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net9209), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net9209), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net9209), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_WIDTH6_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_15 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net9227;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_15 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9227), .TE(1'b0) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net9227), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net9227), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net9227), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net9227), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net9227), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net9227), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net9227), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net9227), .XR(arstz), .Q(rdat[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_15 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_6_00000002 ( clk, arstz, we, wdat, rdat );
  input [5:0] wdat;
  output [5:0] rdat;
  input clk, arstz, we;
  wire   net9245;

  SNPS_CLOCK_GATE_HIGH_glreg_6_00000002 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9245), .TE(1'b0) );
  DFFSQX1 mem_reg_1_ ( .D(wdat[1]), .C(net9245), .XS(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net9245), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net9245), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net9245), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net9245), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net9245), .XR(arstz), .Q(rdat[5]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_6_00000002 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_WIDTH1_2 ( clk, arstz, we, wdat, rdat );
  input [0:0] wdat;
  output [0:0] rdat;
  input clk, arstz, we;
  wire   n2;

  DFFRQX1 mem_reg_0_ ( .D(n2), .C(clk), .XR(arstz), .Q(rdat[0]) );
  AO22AXL U2 ( .A(we), .B(wdat[0]), .C(rdat[0]), .D(we), .Y(n2) );
endmodule


module glreg_a0_16 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net9263;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_16 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9263), .TE(1'b0) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net9263), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net9263), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net9263), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net9263), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net9263), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net9263), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net9263), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net9263), .XR(arstz), .Q(rdat[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_16 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_17 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net9281;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_17 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9281), .TE(1'b0) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net9281), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net9281), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net9281), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net9281), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net9281), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net9281), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net9281), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net9281), .XR(arstz), .Q(rdat[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_17 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_18 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net9299;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_18 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9299), .TE(1'b0) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net9299), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net9299), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net9299), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net9299), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net9299), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net9299), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net9299), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net9299), .XR(arstz), .Q(rdat[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_18 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module cvctl_a0 ( r_cvcwr, wdat, r_sdischg, r_vcomp, r_idacsh, r_cvofsx, 
        r_cvofs, sdischg_duty, r_hlsb_en, r_hlsb_sel, r_hlsb_freq, r_hlsb_duty, 
        r_fw_pwrv, r_dac0, r_dac3, clk_100k, clk, srstz );
  input [5:0] r_cvcwr;
  input [7:0] wdat;
  output [7:0] r_sdischg;
  output [7:0] r_vcomp;
  output [7:0] r_idacsh;
  output [7:0] r_cvofsx;
  output [15:0] r_cvofs;
  input [11:0] r_fw_pwrv;
  output [10:0] r_dac0;
  output [5:0] r_dac3;
  input r_hlsb_en, r_hlsb_sel, r_hlsb_freq, r_hlsb_duty, clk_100k, clk, srstz;
  output sdischg_duty;
  wire   clk_5k, N29, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N46,
         N47, N84, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99,
         N106, N107, N108, N109, N115, N120, N121, N122, N123, N124, N125,
         N126, N127, N128, N129, N130, net9317, n81, N83, N82, N81, N80, N79,
         N78, N77, N76, N75, N74, N73, N72, N68, N67, N66, N65, N64, N63, N62,
         N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48,
         sub_62_carry_2_, sub_62_carry_3_, sub_62_carry_4_, sub_62_carry_5_,
         n1, n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38;
  wire   [4:0] div20_cnt;
  wire   [10:1] cv_code;
  wire   [4:0] sdischg_cnt;
  wire   [4:2] add_81_carry;
  wire   [4:2] add_41_carry;
  wire   [7:1] add_3_root_sub_0_root_add_46_3_carry;

  glreg_a0_24 u0_v_comp ( .clk(clk), .arstz(n8), .we(r_cvcwr[3]), .wdat(wdat), 
        .rdat(r_vcomp) );
  glreg_a0_23 u0_idac_shift ( .clk(clk), .arstz(n7), .we(r_cvcwr[4]), .wdat(
        wdat), .rdat(r_idacsh) );
  glreg_a0_22 u0_cv_ofsx ( .clk(clk), .arstz(n6), .we(r_cvcwr[5]), .wdat(wdat), 
        .rdat(r_cvofsx) );
  glreg_a0_21 u0_cvofs01 ( .clk(clk), .arstz(n5), .we(r_cvcwr[0]), .wdat(wdat), 
        .rdat(r_cvofs[7:0]) );
  glreg_a0_20 u0_cvofs23 ( .clk(clk), .arstz(n4), .we(r_cvcwr[1]), .wdat(wdat), 
        .rdat(r_cvofs[15:8]) );
  glreg_a0_19 u0_sdischg ( .clk(clk), .arstz(n2), .we(r_cvcwr[2]), .wdat(wdat), 
        .rdat(r_sdischg) );
  SNPS_CLOCK_GATE_HIGH_cvctl_a0 clk_gate_sdischg_cnt_reg ( .CLK(clk_100k), 
        .EN(N115), .ENCLK(net9317), .TE(1'b0) );
  cvctl_a0_DW01_add_0 add_62 ( .A({N99, N98, N97, N96, N95, N94}), .B({1'b0, 
        1'b0, N109, N108, N107, N106}), .CI(1'b0), .SUM(r_dac3), .CO() );
  cvctl_a0_DW01_sub_1 sub_2_root_sub_0_root_add_46_3 ( .A(r_fw_pwrv), .B({1'b0, 
        1'b0, 1'b0, 1'b0, r_idacsh}), .CI(1'b0), .DIFF({N59, N58, N57, N56, 
        N55, N54, N53, N52, N51, N50, N49, N48}), .CO() );
  cvctl_a0_DW01_add_2 add_1_root_sub_0_root_add_46_3 ( .A({r_cvofsx[7], 
        r_cvofsx[7], r_cvofsx[7], r_cvofsx[7], r_cvofsx}), .B({1'b0, 1'b0, 
        1'b0, N68, N67, N66, N65, N64, N63, N62, N61, N60}), .CI(1'b0), .SUM({
        N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72}), .CO() );
  cvctl_a0_DW01_add_1 add_0_root_sub_0_root_add_46_3 ( .A({N59, N58, N57, N56, 
        N55, N54, N53, N52, N51, N50, N49, N48}), .B({N83, N82, N81, N80, N79, 
        N78, N77, N76, N75, N74, N73, N72}), .CI(1'b0), .SUM({N84, cv_code, 
        r_dac0[0]}), .CO() );
  HAD1X1 add_81_U1_1_1 ( .A(sdischg_cnt[1]), .B(sdischg_cnt[0]), .CO(
        add_81_carry[2]), .SO(N121) );
  HAD1X1 add_81_U1_1_2 ( .A(sdischg_cnt[2]), .B(add_81_carry[2]), .CO(
        add_81_carry[3]), .SO(N122) );
  HAD1X1 add_81_U1_1_3 ( .A(sdischg_cnt[3]), .B(add_81_carry[3]), .CO(
        add_81_carry[4]), .SO(N123) );
  HAD1X1 add_41_U1_1_1 ( .A(div20_cnt[1]), .B(div20_cnt[0]), .CO(
        add_41_carry[2]), .SO(N34) );
  HAD1X1 add_41_U1_1_2 ( .A(div20_cnt[2]), .B(add_41_carry[2]), .CO(
        add_41_carry[3]), .SO(N35) );
  HAD1X1 add_41_U1_1_3 ( .A(div20_cnt[3]), .B(add_41_carry[3]), .CO(
        add_41_carry[4]), .SO(N36) );
  FAD1X1 add_3_root_sub_0_root_add_46_3_U1_1 ( .A(N47), .B(r_vcomp[1]), .CI(
        add_3_root_sub_0_root_add_46_3_carry[1]), .CO(
        add_3_root_sub_0_root_add_46_3_carry[2]), .SO(N61) );
  DFFRQX1 sdischg_cnt_reg_4_ ( .D(N130), .C(net9317), .XR(n6), .Q(
        sdischg_cnt[4]) );
  DFFRQX1 sdischg_cnt_reg_0_ ( .D(N126), .C(net9317), .XR(srstz), .Q(
        sdischg_cnt[0]) );
  DFFRQX1 div20_cnt_reg_1_ ( .D(N39), .C(clk_100k), .XR(n5), .Q(div20_cnt[1])
         );
  DFFRQX1 div20_cnt_reg_3_ ( .D(N41), .C(clk_100k), .XR(n4), .Q(div20_cnt[3])
         );
  DFFRQX1 div20_cnt_reg_0_ ( .D(N38), .C(clk_100k), .XR(n8), .Q(div20_cnt[0])
         );
  DFFRQX1 div20_cnt_reg_2_ ( .D(N40), .C(clk_100k), .XR(n2), .Q(div20_cnt[2])
         );
  DFFRQX1 div20_cnt_reg_4_ ( .D(N42), .C(clk_100k), .XR(n8), .Q(div20_cnt[4])
         );
  DFFRQX1 sdischg_cnt_reg_2_ ( .D(N128), .C(net9317), .XR(n4), .Q(
        sdischg_cnt[2]) );
  DFFRQX1 sdischg_cnt_reg_3_ ( .D(N129), .C(net9317), .XR(n7), .Q(
        sdischg_cnt[3]) );
  DFFRQX1 sdischg_cnt_reg_1_ ( .D(N127), .C(net9317), .XR(srstz), .Q(
        sdischg_cnt[1]) );
  DFFRQX1 sdischg_reg ( .D(n81), .C(net9317), .XR(n6), .Q(sdischg_duty) );
  DFFRQX1 clk_5k_reg ( .D(N29), .C(clk_100k), .XR(n5), .Q(clk_5k) );
  INVX1 U3 ( .A(n37), .Y(n1) );
  INVX1 U4 ( .A(n9), .Y(n8) );
  INVX1 U5 ( .A(n9), .Y(n4) );
  INVX1 U6 ( .A(n9), .Y(n5) );
  INVX1 U7 ( .A(n9), .Y(n6) );
  INVX1 U8 ( .A(n9), .Y(n7) );
  INVX1 U9 ( .A(n9), .Y(n2) );
  INVX1 U10 ( .A(srstz), .Y(n9) );
  INVX1 U12 ( .A(r_sdischg[3]), .Y(n18) );
  INVX1 U13 ( .A(sdischg_cnt[1]), .Y(n16) );
  INVX1 U14 ( .A(r_sdischg[2]), .Y(n17) );
  INVX1 U15 ( .A(r_sdischg[4]), .Y(n19) );
  AND2X1 U16 ( .A(r_vcomp[7]), .B(add_3_root_sub_0_root_add_46_3_carry[7]), 
        .Y(N68) );
  XOR2X1 U17 ( .A(add_3_root_sub_0_root_add_46_3_carry[7]), .B(r_vcomp[7]), 
        .Y(N67) );
  XOR2X1 U18 ( .A(cv_code[6]), .B(sub_62_carry_5_), .Y(N93) );
  AND2X1 U19 ( .A(cv_code[5]), .B(sub_62_carry_4_), .Y(sub_62_carry_5_) );
  XOR2X1 U20 ( .A(sub_62_carry_4_), .B(cv_code[5]), .Y(N92) );
  AND2X1 U21 ( .A(cv_code[4]), .B(sub_62_carry_3_), .Y(sub_62_carry_4_) );
  XOR2X1 U22 ( .A(sub_62_carry_3_), .B(cv_code[4]), .Y(N91) );
  AND2X1 U23 ( .A(cv_code[3]), .B(sub_62_carry_2_), .Y(sub_62_carry_3_) );
  XOR2X1 U24 ( .A(sub_62_carry_2_), .B(cv_code[3]), .Y(N90) );
  AND2X1 U25 ( .A(cv_code[2]), .B(cv_code[1]), .Y(sub_62_carry_2_) );
  XOR2X1 U26 ( .A(cv_code[1]), .B(cv_code[2]), .Y(N89) );
  AND2X1 U27 ( .A(r_vcomp[6]), .B(add_3_root_sub_0_root_add_46_3_carry[6]), 
        .Y(add_3_root_sub_0_root_add_46_3_carry[7]) );
  XOR2X1 U28 ( .A(add_3_root_sub_0_root_add_46_3_carry[6]), .B(r_vcomp[6]), 
        .Y(N66) );
  AND2X1 U29 ( .A(r_vcomp[5]), .B(add_3_root_sub_0_root_add_46_3_carry[5]), 
        .Y(add_3_root_sub_0_root_add_46_3_carry[6]) );
  XOR2X1 U30 ( .A(add_3_root_sub_0_root_add_46_3_carry[5]), .B(r_vcomp[5]), 
        .Y(N65) );
  AND2X1 U31 ( .A(r_vcomp[4]), .B(add_3_root_sub_0_root_add_46_3_carry[4]), 
        .Y(add_3_root_sub_0_root_add_46_3_carry[5]) );
  XOR2X1 U32 ( .A(add_3_root_sub_0_root_add_46_3_carry[4]), .B(r_vcomp[4]), 
        .Y(N64) );
  AND2X1 U33 ( .A(r_vcomp[3]), .B(add_3_root_sub_0_root_add_46_3_carry[3]), 
        .Y(add_3_root_sub_0_root_add_46_3_carry[4]) );
  XOR2X1 U34 ( .A(add_3_root_sub_0_root_add_46_3_carry[3]), .B(r_vcomp[3]), 
        .Y(N63) );
  AND2X1 U35 ( .A(r_vcomp[2]), .B(add_3_root_sub_0_root_add_46_3_carry[2]), 
        .Y(add_3_root_sub_0_root_add_46_3_carry[3]) );
  XOR2X1 U36 ( .A(add_3_root_sub_0_root_add_46_3_carry[2]), .B(r_vcomp[2]), 
        .Y(N62) );
  AND2X1 U37 ( .A(r_vcomp[0]), .B(N46), .Y(
        add_3_root_sub_0_root_add_46_3_carry[1]) );
  XOR2X1 U38 ( .A(N46), .B(r_vcomp[0]), .Y(N60) );
  INVX1 U39 ( .A(cv_code[1]), .Y(N88) );
  INVX1 U40 ( .A(div20_cnt[0]), .Y(N33) );
  XOR2X1 U41 ( .A(add_41_carry[4]), .B(div20_cnt[4]), .Y(N37) );
  INVX1 U42 ( .A(sdischg_cnt[0]), .Y(N120) );
  XOR2X1 U43 ( .A(add_81_carry[4]), .B(sdischg_cnt[4]), .Y(N124) );
  AND2X1 U44 ( .A(sdischg_cnt[3]), .B(n18), .Y(n11) );
  OAI32X1 U45 ( .A(n17), .B(sdischg_cnt[2]), .C(n11), .D(sdischg_cnt[3]), .E(
        n18), .Y(n12) );
  AOI22BXL U46 ( .B(r_sdischg[1]), .A(sdischg_cnt[1]), .D(r_sdischg[0]), .C(
        sdischg_cnt[0]), .Y(n10) );
  AOI211X1 U47 ( .C(r_sdischg[1]), .D(n16), .A(n12), .B(n10), .Y(n15) );
  AOI21X1 U48 ( .B(sdischg_cnt[2]), .C(n17), .A(n11), .Y(n13) );
  ENOX1 U49 ( .A(n13), .B(n12), .C(n19), .D(sdischg_cnt[4]), .Y(n14) );
  OAI22X1 U50 ( .A(sdischg_cnt[4]), .B(n19), .C(n15), .D(n14), .Y(N125) );
  OR2X1 U51 ( .A(cv_code[8]), .B(n1), .Y(r_dac0[8]) );
  OR2X1 U52 ( .A(cv_code[7]), .B(n1), .Y(r_dac0[7]) );
  OR2X1 U53 ( .A(cv_code[6]), .B(n1), .Y(r_dac0[6]) );
  OR2X1 U54 ( .A(cv_code[5]), .B(n1), .Y(r_dac0[5]) );
  OR2X1 U55 ( .A(cv_code[4]), .B(n1), .Y(r_dac0[4]) );
  OR2X1 U56 ( .A(cv_code[3]), .B(n1), .Y(r_dac0[3]) );
  OR2X1 U57 ( .A(cv_code[2]), .B(N84), .Y(r_dac0[2]) );
  OR2X1 U58 ( .A(cv_code[1]), .B(N84), .Y(r_dac0[1]) );
  MUX2X1 U59 ( .D0(N125), .D1(sdischg_duty), .S(n20), .Y(n81) );
  AND2X1 U60 ( .A(N93), .B(N84), .Y(N99) );
  AND2X1 U61 ( .A(N92), .B(N84), .Y(N98) );
  AND2X1 U62 ( .A(N91), .B(N84), .Y(N97) );
  AND2X1 U63 ( .A(N90), .B(N84), .Y(N96) );
  AND2X1 U64 ( .A(N89), .B(N84), .Y(N95) );
  AND2X1 U65 ( .A(N88), .B(N84), .Y(N94) );
  NOR32XL U66 ( .B(r_hlsb_en), .C(clk_5k), .A(r_hlsb_sel), .Y(N47) );
  NOR32XL U67 ( .B(r_hlsb_sel), .C(clk_5k), .A(n21), .Y(N46) );
  NOR21XL U68 ( .B(N37), .A(n22), .Y(N42) );
  NOR21XL U69 ( .B(N36), .A(n22), .Y(N41) );
  NOR21XL U70 ( .B(N35), .A(n22), .Y(N40) );
  NOR21XL U71 ( .B(N34), .A(n22), .Y(N39) );
  NOR21XL U72 ( .B(N33), .A(n22), .Y(N38) );
  OAI221X1 U73 ( .A(n23), .B(n24), .C(n25), .D(n26), .E(r_hlsb_en), .Y(n22) );
  AOI221XL U74 ( .A(div20_cnt[3]), .B(n24), .C(div20_cnt[1]), .D(div20_cnt[0]), 
        .E(div20_cnt[2]), .Y(n25) );
  INVX1 U75 ( .A(r_hlsb_freq), .Y(n24) );
  AOI21BX1 U76 ( .C(n26), .B(n27), .A(div20_cnt[4]), .Y(n23) );
  MUX2IX1 U77 ( .D0(div20_cnt[4]), .D1(div20_cnt[3]), .S(r_hlsb_freq), .Y(n26)
         );
  AOI31X1 U78 ( .A(n28), .B(n29), .C(n30), .D(n21), .Y(N29) );
  INVX1 U79 ( .A(r_hlsb_en), .Y(n21) );
  OAI31XL U80 ( .A(n31), .B(r_hlsb_freq), .C(div20_cnt[2]), .D(div20_cnt[3]), 
        .Y(n30) );
  AO21X1 U81 ( .B(div20_cnt[0]), .C(r_hlsb_duty), .A(div20_cnt[1]), .Y(n31) );
  INVX1 U82 ( .A(div20_cnt[4]), .Y(n29) );
  OAI211X1 U83 ( .C(r_hlsb_duty), .D(n27), .A(r_hlsb_freq), .B(div20_cnt[2]), 
        .Y(n28) );
  OR2X1 U84 ( .A(div20_cnt[0]), .B(div20_cnt[1]), .Y(n27) );
  NOR21XL U85 ( .B(N124), .A(n20), .Y(N130) );
  NOR21XL U86 ( .B(N123), .A(n20), .Y(N129) );
  NOR21XL U87 ( .B(N122), .A(n20), .Y(N128) );
  NOR21XL U88 ( .B(N121), .A(n20), .Y(N127) );
  NOR21XL U89 ( .B(N120), .A(n20), .Y(N126) );
  NAND42X1 U90 ( .C(sdischg_cnt[1]), .D(sdischg_cnt[0]), .A(n20), .B(n32), .Y(
        N115) );
  NOR3XL U91 ( .A(sdischg_cnt[2]), .B(sdischg_cnt[4]), .C(sdischg_cnt[3]), .Y(
        n32) );
  NOR2X1 U92 ( .A(r_sdischg[6]), .B(r_sdischg[5]), .Y(n20) );
  AO2222XL U93 ( .A(r_cvofs[7]), .B(n33), .C(r_cvofs[15]), .D(n34), .E(
        r_cvofs[14]), .F(n35), .G(r_cvofs[6]), .H(n36), .Y(N109) );
  AO2222XL U94 ( .A(r_cvofs[2]), .B(n33), .C(r_cvofs[10]), .D(n34), .E(
        r_cvofs[13]), .F(n35), .G(r_cvofs[5]), .H(n36), .Y(N108) );
  AO2222XL U95 ( .A(r_cvofs[1]), .B(n33), .C(r_cvofs[9]), .D(n34), .E(
        r_cvofs[12]), .F(n35), .G(r_cvofs[4]), .H(n36), .Y(N107) );
  AO2222XL U96 ( .A(r_cvofs[0]), .B(n33), .C(r_cvofs[8]), .D(n34), .E(
        r_cvofs[11]), .F(n35), .G(r_cvofs[3]), .H(n36), .Y(N106) );
  NOR2X1 U97 ( .A(n33), .B(r_dac0[10]), .Y(n36) );
  OAI21BBX1 U98 ( .A(cv_code[10]), .B(cv_code[9]), .C(n37), .Y(n35) );
  NOR2X1 U99 ( .A(n38), .B(r_dac0[9]), .Y(n34) );
  NAND21X1 U100 ( .B(cv_code[9]), .A(n37), .Y(r_dac0[9]) );
  INVX1 U101 ( .A(N84), .Y(n37) );
  NOR2X1 U102 ( .A(r_dac0[10]), .B(cv_code[9]), .Y(n33) );
  INVX1 U103 ( .A(n38), .Y(r_dac0[10]) );
  NOR2X1 U104 ( .A(cv_code[10]), .B(N84), .Y(n38) );
endmodule


module cvctl_a0_DW01_add_1 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;

  wire   [11:1] carry;

  FAD1X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .SO(
        SUM[10]) );
  FAD1X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .SO(SUM[9])
         );
  FAD1X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .SO(SUM[8])
         );
  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  XOR3X1 U1_11 ( .A(A[11]), .B(B[11]), .C(carry[11]), .Y(SUM[11]) );
  AND2X1 U1 ( .A(A[0]), .B(B[0]), .Y(carry[1]) );
  XOR2X1 U2 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
endmodule


module cvctl_a0_DW01_add_2 ( A, B, CI, SUM, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;

  wire   [11:1] carry;

  FAD1X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .SO(SUM[8])
         );
  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  XOR2X1 U1 ( .A(carry[9]), .B(A[9]), .Y(SUM[9]) );
  XOR2X1 U2 ( .A(carry[10]), .B(A[10]), .Y(SUM[10]) );
  XOR2X1 U3 ( .A(A[11]), .B(carry[11]), .Y(SUM[11]) );
  AND2X1 U4 ( .A(A[0]), .B(B[0]), .Y(carry[1]) );
  XOR2X1 U5 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
  AND2X1 U6 ( .A(carry[9]), .B(A[9]), .Y(carry[10]) );
  AND2X1 U7 ( .A(carry[10]), .B(A[10]), .Y(carry[11]) );
endmodule


module cvctl_a0_DW01_sub_1 ( A, B, CI, DIFF, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10;
  wire   [10:1] carry;

  FAD1X1 U2_7 ( .A(A[7]), .B(n3), .CI(carry[7]), .CO(carry[8]), .SO(DIFF[7])
         );
  FAD1X1 U2_6 ( .A(A[6]), .B(n4), .CI(carry[6]), .CO(carry[7]), .SO(DIFF[6])
         );
  FAD1X1 U2_5 ( .A(A[5]), .B(n5), .CI(carry[5]), .CO(carry[6]), .SO(DIFF[5])
         );
  FAD1X1 U2_4 ( .A(A[4]), .B(n6), .CI(carry[4]), .CO(carry[5]), .SO(DIFF[4])
         );
  FAD1X1 U2_3 ( .A(A[3]), .B(n7), .CI(carry[3]), .CO(carry[4]), .SO(DIFF[3])
         );
  FAD1X1 U2_2 ( .A(A[2]), .B(n8), .CI(carry[2]), .CO(carry[3]), .SO(DIFF[2])
         );
  FAD1X1 U2_1 ( .A(A[1]), .B(n9), .CI(carry[1]), .CO(carry[2]), .SO(DIFF[1])
         );
  NOR2X1 U1 ( .A(A[10]), .B(carry[10]), .Y(n1) );
  XOR2X1 U2 ( .A(n1), .B(A[11]), .Y(DIFF[11]) );
  XNOR2XL U3 ( .A(A[8]), .B(carry[8]), .Y(DIFF[8]) );
  XNOR2XL U4 ( .A(A[9]), .B(carry[9]), .Y(DIFF[9]) );
  XNOR2XL U5 ( .A(A[10]), .B(carry[10]), .Y(DIFF[10]) );
  INVX1 U6 ( .A(B[7]), .Y(n3) );
  INVX1 U7 ( .A(B[2]), .Y(n8) );
  INVX1 U8 ( .A(B[3]), .Y(n7) );
  INVX1 U9 ( .A(B[4]), .Y(n6) );
  INVX1 U10 ( .A(B[5]), .Y(n5) );
  INVX1 U11 ( .A(B[6]), .Y(n4) );
  INVX1 U12 ( .A(B[1]), .Y(n9) );
  NAND21X1 U13 ( .B(n10), .A(n2), .Y(carry[1]) );
  INVX1 U14 ( .A(A[0]), .Y(n2) );
  OR2X1 U15 ( .A(A[8]), .B(carry[8]), .Y(carry[9]) );
  XNOR2XL U16 ( .A(n10), .B(A[0]), .Y(DIFF[0]) );
  INVX1 U17 ( .A(B[0]), .Y(n10) );
  OR2X1 U18 ( .A(A[9]), .B(carry[9]), .Y(carry[10]) );
endmodule


module cvctl_a0_DW01_add_0 ( A, B, CI, SUM, CO );
  input [5:0] A;
  input [5:0] B;
  output [5:0] SUM;
  input CI;
  output CO;
  wire   n1, n2;
  wire   [5:1] carry;

  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  INVX1 U1 ( .A(A[4]), .Y(n1) );
  INVX1 U2 ( .A(B[0]), .Y(n2) );
  XOR2X1 U3 ( .A(A[5]), .B(carry[5]), .Y(SUM[5]) );
  NOR21XL U4 ( .B(carry[4]), .A(n1), .Y(carry[5]) );
  XOR2X1 U5 ( .A(carry[4]), .B(A[4]), .Y(SUM[4]) );
  XOR2X1 U6 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
  NOR21XL U7 ( .B(A[0]), .A(n2), .Y(carry[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_cvctl_a0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_19 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net9335;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_19 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9335), .TE(1'b0) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net9335), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net9335), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net9335), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net9335), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net9335), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net9335), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net9335), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net9335), .XR(arstz), .Q(rdat[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_19 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_20 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net9353;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_20 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9353), .TE(1'b0) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net9353), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net9353), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net9353), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net9353), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net9353), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net9353), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net9353), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net9353), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_20 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_21 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net9371;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_21 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9371), .TE(1'b0) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net9371), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net9371), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net9371), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net9371), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net9371), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net9371), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net9371), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net9371), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_21 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_22 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net9389;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_22 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9389), .TE(1'b0) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net9389), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net9389), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net9389), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net9389), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net9389), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net9389), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net9389), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net9389), .XR(arstz), .Q(rdat[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_22 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_23 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net9407;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_23 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9407), .TE(1'b0) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net9407), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net9407), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net9407), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net9407), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net9407), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net9407), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net9407), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net9407), .XR(arstz), .Q(rdat[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_23 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_24 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net9425;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_24 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9425), .TE(1'b0) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net9425), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net9425), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net9425), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net9425), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net9425), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net9425), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net9425), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net9425), .XR(arstz), .Q(rdat[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_24 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module fcp_a0 ( dp_comp, dm_comp, id_comp, intr, tx_en, tx_dat, r_dat, r_sta, 
        r_ctl, r_msk, r_crc, r_acc, r_dpdmsta, r_wdat, r_wr, r_re, clk, srstz, 
        r_tui );
  output [7:0] r_dat;
  output [7:0] r_sta;
  output [7:0] r_ctl;
  output [7:0] r_msk;
  output [7:0] r_crc;
  output [7:0] r_acc;
  output [7:0] r_dpdmsta;
  input [7:0] r_wdat;
  input [6:0] r_wr;
  output [7:0] r_tui;
  input dp_comp, dm_comp, id_comp, r_re, clk, srstz;
  output intr, tx_en, tx_dat;
  wire   r_dm, r_dmchg, r_acc_int, r_wr_last, r_wr_other, n1, n2, n3, n4;

  dpdmacc_a0 u0_dpdmacc ( .dp_comp(dp_comp), .dm_comp(dm_comp), .id_comp(
        id_comp), .r_re_0(r_re), .r_wr_1(r_wr[6]), .r_wdat(r_wdat), .r_acc(
        r_acc), .r_dpdmsta(r_dpdmsta), .r_dm(r_dm), .r_dmchg(r_dmchg), .r_int(
        r_acc_int), .clk(clk), .rstz(srstz) );
  fcpegn_a0 u0_fcpegn ( .intr(intr), .tx_en(tx_en), .tx_dat(tx_dat), .r_dat(
        r_dat), .r_sta(r_sta), .r_ctl(r_ctl), .r_msk(r_msk), .r_wr(r_wr[4:0]), 
        .r_wdat(r_wdat), .ff_idn(n2), .ff_chg(n1), .r_acc_int(r_acc_int), 
        .clk(clk), .srstz(n3), .r_tui(r_tui) );
  fcpcrc_a0 u0_fcpcrc ( .tx_crc(r_crc), .crc_din(r_wdat), .crc_en(r_ctl[2]), 
        .crc_shfi(r_wr_other), .crc_shfl(r_wr_last), .clk(clk), .srstz(n3) );
  BUFX3 U1 ( .A(r_dmchg), .Y(n1) );
  BUFX3 U2 ( .A(r_dm), .Y(n2) );
  INVX1 U3 ( .A(n4), .Y(n3) );
  INVX1 U4 ( .A(srstz), .Y(n4) );
  AND2X1 U5 ( .A(r_wr[5]), .B(r_ctl[3]), .Y(r_wr_last) );
  NOR21XL U6 ( .B(r_wr[5]), .A(r_ctl[3]), .Y(r_wr_other) );
endmodule


module fcpcrc_a0 ( tx_crc, crc_din, crc_en, crc_shfi, crc_shfl, clk, srstz );
  output [7:0] tx_crc;
  input [7:0] crc_din;
  input crc_en, crc_shfi, crc_shfl, clk, srstz;
  wire   N81, N82, N83, N84, N85, N86, N87, N88, N89, net9443, n3, n4, n5, n6,
         n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n1, n2;

  SNPS_CLOCK_GATE_HIGH_fcpcrc_a0 clk_gate_crc8_r_reg ( .CLK(clk), .EN(N81), 
        .ENCLK(net9443), .TE(1'b0) );
  DFFRQX1 crc8_r_reg_2_ ( .D(N84), .C(net9443), .XR(srstz), .Q(tx_crc[2]) );
  DFFRQX1 crc8_r_reg_0_ ( .D(N82), .C(net9443), .XR(srstz), .Q(tx_crc[0]) );
  DFFRQX1 crc8_r_reg_3_ ( .D(N85), .C(net9443), .XR(srstz), .Q(tx_crc[3]) );
  DFFRQX1 crc8_r_reg_1_ ( .D(N83), .C(net9443), .XR(srstz), .Q(tx_crc[1]) );
  DFFRQX1 crc8_r_reg_6_ ( .D(N88), .C(net9443), .XR(srstz), .Q(tx_crc[6]) );
  DFFRQX1 crc8_r_reg_7_ ( .D(N89), .C(net9443), .XR(srstz), .Q(tx_crc[7]) );
  DFFRQX1 crc8_r_reg_5_ ( .D(N87), .C(net9443), .XR(srstz), .Q(tx_crc[5]) );
  DFFRQX1 crc8_r_reg_4_ ( .D(N86), .C(net9443), .XR(srstz), .Q(tx_crc[4]) );
  XNOR2XL U3 ( .A(n29), .B(n26), .Y(n15) );
  XNOR2XL U4 ( .A(n15), .B(n24), .Y(n8) );
  XNOR2XL U5 ( .A(n35), .B(n34), .Y(n20) );
  XNOR2XL U6 ( .A(n8), .B(n17), .Y(n35) );
  XNOR2XL U7 ( .A(n28), .B(n29), .Y(n9) );
  XNOR2XL U8 ( .A(n17), .B(n27), .Y(n28) );
  XNOR2XL U9 ( .A(crc_din[1]), .B(n1), .Y(n31) );
  XNOR2XL U10 ( .A(n5), .B(n11), .Y(n29) );
  OAI22X1 U11 ( .A(n16), .B(n4), .C(n17), .D(n6), .Y(N87) );
  XNOR2XL U12 ( .A(n18), .B(n19), .Y(n16) );
  XNOR2XL U13 ( .A(n9), .B(n17), .Y(n19) );
  XNOR2XL U14 ( .A(n20), .B(n14), .Y(n18) );
  OAI22X1 U15 ( .A(n4), .B(n21), .C(n22), .D(n6), .Y(N86) );
  XOR2X1 U16 ( .A(n20), .B(n23), .Y(n21) );
  XOR2X1 U17 ( .A(n14), .B(n24), .Y(n23) );
  OAI22X1 U18 ( .A(n25), .B(n4), .C(n26), .D(n6), .Y(N85) );
  XNOR2XL U19 ( .A(n20), .B(n15), .Y(n25) );
  OAI22X1 U20 ( .A(n4), .B(n20), .C(n34), .D(n6), .Y(N82) );
  XNOR2XL U21 ( .A(n37), .B(n38), .Y(n17) );
  XNOR2XL U22 ( .A(n30), .B(n39), .Y(n38) );
  XNOR2XL U23 ( .A(crc_din[5]), .B(n2), .Y(n39) );
  XNOR2XL U24 ( .A(n32), .B(n33), .Y(n14) );
  XNOR2XL U25 ( .A(n17), .B(n11), .Y(n33) );
  XNOR2XL U26 ( .A(n24), .B(n31), .Y(n32) );
  XNOR2XL U27 ( .A(n22), .B(n5), .Y(n24) );
  XNOR2XL U28 ( .A(n37), .B(n40), .Y(n22) );
  XOR2X1 U29 ( .A(crc_din[4]), .B(n41), .Y(n40) );
  XNOR2XL U30 ( .A(n36), .B(n43), .Y(n26) );
  XOR2X1 U31 ( .A(crc_din[3]), .B(n44), .Y(n43) );
  OAI22X1 U32 ( .A(n10), .B(n4), .C(n11), .D(n6), .Y(N88) );
  XNOR2XL U33 ( .A(n12), .B(n13), .Y(n10) );
  XNOR2XL U34 ( .A(n14), .B(n15), .Y(n12) );
  XNOR2XL U35 ( .A(n9), .B(n11), .Y(n13) );
  OAI22X1 U36 ( .A(n3), .B(n4), .C(n5), .D(n6), .Y(N89) );
  XNOR2XL U37 ( .A(n7), .B(n8), .Y(n3) );
  XNOR2XL U38 ( .A(n9), .B(n5), .Y(n7) );
  OAI22X1 U39 ( .A(n4), .B(n14), .C(n31), .D(n6), .Y(N83) );
  OAI22X1 U40 ( .A(n9), .B(n4), .C(n27), .D(n6), .Y(N84) );
  XNOR2XL U41 ( .A(crc_din[2]), .B(n30), .Y(n27) );
  XNOR2XL U42 ( .A(crc_din[0]), .B(n36), .Y(n34) );
  XNOR2XL U43 ( .A(n36), .B(n1), .Y(n37) );
  XNOR2XL U44 ( .A(n44), .B(n41), .Y(n45) );
  INVX1 U45 ( .A(n42), .Y(n1) );
  XNOR2XL U46 ( .A(n47), .B(n48), .Y(n11) );
  XNOR2XL U47 ( .A(n42), .B(n30), .Y(n48) );
  XNOR2XL U48 ( .A(n44), .B(n51), .Y(n47) );
  XNOR2XL U49 ( .A(tx_crc[6]), .B(crc_din[6]), .Y(n51) );
  XNOR2XL U50 ( .A(n52), .B(n53), .Y(n5) );
  XNOR2XL U51 ( .A(n45), .B(n30), .Y(n52) );
  XNOR2XL U52 ( .A(tx_crc[7]), .B(crc_din[7]), .Y(n53) );
  NAND21X1 U53 ( .B(crc_shfl), .A(crc_en), .Y(n6) );
  NAND2X1 U54 ( .A(crc_shfl), .B(crc_en), .Y(n4) );
  OR2X1 U55 ( .A(crc_shfi), .B(n6), .Y(N81) );
  XNOR2XL U56 ( .A(n49), .B(n50), .Y(n42) );
  XNOR2XL U57 ( .A(n2), .B(tx_crc[6]), .Y(n49) );
  XNOR2XL U58 ( .A(tx_crc[1]), .B(n41), .Y(n50) );
  XOR2X1 U59 ( .A(n54), .B(n55), .Y(n30) );
  XNOR2XL U60 ( .A(tx_crc[5]), .B(tx_crc[2]), .Y(n54) );
  XOR2X1 U61 ( .A(n45), .B(n46), .Y(n36) );
  XNOR2XL U62 ( .A(tx_crc[0]), .B(n2), .Y(n46) );
  XNOR2XL U63 ( .A(tx_crc[3]), .B(n55), .Y(n44) );
  XNOR2XL U64 ( .A(tx_crc[7]), .B(tx_crc[4]), .Y(n41) );
  XNOR2XL U65 ( .A(tx_crc[7]), .B(tx_crc[6]), .Y(n55) );
  INVX1 U66 ( .A(tx_crc[5]), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_fcpcrc_a0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module fcpegn_a0 ( intr, tx_en, tx_dat, r_dat, r_sta, r_ctl, r_msk, r_wr, 
        r_wdat, ff_idn, ff_chg, r_acc_int, clk, srstz, r_tui );
  output [7:0] r_dat;
  output [7:0] r_sta;
  output [7:0] r_ctl;
  output [7:0] r_msk;
  input [4:0] r_wr;
  input [7:0] r_wdat;
  output [7:0] r_tui;
  input ff_idn, ff_chg, r_acc_int, clk, srstz;
  output intr, tx_en, tx_dat;
  wire   N22, upd_dbuf_en, N85, N87, N88, N95, N96, N97, N98, N99, N141, N142,
         N143, N144, N145, N146, N147, N148, N149, N150, N151, N152, N153,
         N171, N172, N173, N174, N175, N176, N177, N178, N179, N180, N181,
         N186, N187, N188, N189, N190, N192, adp_tx_ui_7_, adp_tx_ui_6_,
         adp_tx_ui_5_, tui_upd, N205, N219, N221, N222, N223, N224, N225, N226,
         N227, N228, N260, N261, N324, N325, N326, N328, N331, N336, N337,
         N338, N348, N349, N356, N362, N363, N418, N419, N444, rx_trans_8_chg,
         N1005, N1006, N1007, N1008, N1009, N1010, N1011, N1012, N1013, N1014,
         N1015, N1016, N1043, net9465, net9469, net9472, net9473, net9474,
         net9475, net9476, net9477, net9480, net9483, net9488, net9493,
         net9498, n26, n27, n28, n29, n30, n31, n32, n516, n517, n525, n526,
         N1259, N1258, N1257, N1256, N1255, N1254, N1253, N1252, N168, N167,
         N166, N165, N164, N163, N162, N161, N160, N159, N116, N115, N114,
         N113, N112, N111, N110, N109, N108, N107, gt_647_B_3_,
         add_423_carry_5_, sub_423_carry_5_, add_264_A_0_, add_282_carry_7_,
         mult_274_2_n7, mult_274_2_n6, mult_274_2_n5, mult_274_2_n4,
         mult_274_2_n3, mult_274_2_n2, mult_274_n7, mult_274_n6, mult_274_n5,
         mult_274_n4, mult_274_n3, mult_274_n2, n1, n2, n3, n4, n5, n6, n7, n8,
         n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n22, n23, n24,
         n25, n33, n34, n35, n36, n37, n38, n39, n40, n41, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461,
         SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2,
         SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4;
  wire   [6:0] setsta;
  wire   [7:0] clrsta;
  wire   [7:0] r_irq;
  wire   [7:0] upd_dbuf;
  wire   [10:0] rxtx_buf;
  wire   [3:0] us_cnt;
  wire   [6:4] rx_ui_1_2;
  wire   [6:0] rx_ui_3_8;
  wire   [7:0] rx_ui_5_8;
  wire   [5:0] catch_sync;
  wire   [7:0] ui_intv_cnt;
  wire   [6:2] symb_cnt;
  wire   [15:3] catch_ping;
  wire   [12:5] ui_by_ping;
  wire   [6:0] adp_tx_1_4;
  wire   [7:0] tui_wdat;
  wire   [11:0] trans_buf;
  wire   [1:0] new_rx_sync_cnt;
  wire   [3:0] fcp_state;
  wire   [11:1] add_277_carry;
  wire   [6:1] add_264_carry;
  wire   [5:1] add_263_carry;
  wire   [14:6] add_274_2_carry;
  wire   [15:6] add_274_carry;

  glreg_8_00000000 u0_fcpctl ( .clk(clk), .arstz(n46), .we(r_wr[0]), .wdat({
        n39, n37, r_wdat[5:3], n25, r_wdat[1:0]}), .rdat({
        SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3, 
        r_ctl[4:0]}) );
  glsta_a0_0 u0_fcpsta ( .clk(clk), .arstz(n45), .rst0(1'b0), .set2({r_acc_int, 
        setsta[6:3], n525, n517, setsta[0]}), .clr1(clrsta), .rdat(r_sta), 
        .irq(r_irq) );
  glreg_a0_4 u0_fcpmsk ( .clk(clk), .arstz(n44), .we(r_wr[2]), .wdat({n39, n37, 
        r_wdat[5:3], n25, r_wdat[1:0]}), .rdat(r_msk) );
  glreg_a0_3 u0_fcpdat ( .clk(clk), .arstz(n43), .we(upd_dbuf_en), .wdat(
        upd_dbuf), .rdat(r_dat) );
  glreg_a0_2 u0_fcptui ( .clk(clk), .arstz(n41), .we(tui_upd), .wdat(tui_wdat), 
        .rdat(r_tui) );
  SNPS_CLOCK_GATE_HIGH_fcpegn_a0_0 clk_gate_catch_sync_reg ( .CLK(clk), .EN(
        n526), .ENCLK(net9465), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_fcpegn_a0_4 clk_gate_ui_intv_cnt_reg ( .CLK(clk), .EN(
        N205), .ENCLK(net9483), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_fcpegn_a0_3 clk_gate_rxtx_buf_reg ( .CLK(clk), .EN(N22), 
        .ENCLK(net9488), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_fcpegn_a0_2 clk_gate_fcp_state_reg ( .CLK(clk), .EN(
        N1005), .ENCLK(net9493), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_fcpegn_a0_1 clk_gate_symb_cnt_reg ( .CLK(clk), .EN(
        N1043), .ENCLK(net9498), .TE(1'b0) );
  fcpegn_a0_DW01_inc_0 r611 ( .A({symb_cnt[6:4], n11, symb_cnt[2], n4, n18}), 
        .SUM({n26, n27, n28, n29, n30, n31, n32}) );
  fcpegn_a0_DW01_inc_1 add_283_round ( .A({1'b0, adp_tx_ui_7_, adp_tx_ui_6_, 
        adp_tx_ui_5_, r_tui[4:1]}), .SUM({adp_tx_1_4, SYNOPSYS_UNCONNECTED_4})
         );
  fcpegn_a0_DW01_inc_2 add_316_aco ( .A({N1259, N1258, N1257, N1256, N1255, 
        N1254, N1253, N1252}), .SUM({N228, N227, N226, N225, N224, N223, N222, 
        N221}) );
  FAD1X1 add_264_U1_1 ( .A(N324), .B(n10), .CI(add_264_carry[1]), .CO(
        add_264_carry[2]), .SO(rx_ui_5_8[1]) );
  FAD1X1 add_264_U1_2 ( .A(N325), .B(rx_ui_1_2[4]), .CI(add_264_carry[2]), 
        .CO(add_264_carry[3]), .SO(rx_ui_5_8[2]) );
  FAD1X1 add_264_U1_3 ( .A(n10), .B(gt_647_B_3_), .CI(add_264_carry[3]), .CO(
        add_264_carry[4]), .SO(rx_ui_5_8[3]) );
  FAD1X1 add_264_U1_4 ( .A(n231), .B(rx_ui_1_2[6]), .CI(add_264_carry[4]), 
        .CO(add_264_carry[5]), .SO(rx_ui_5_8[4]) );
  FAD1X1 add_263_U1_1 ( .A(N325), .B(n9), .CI(add_263_carry[1]), .CO(
        add_263_carry[2]), .SO(rx_ui_3_8[1]) );
  FAD1X1 add_263_U1_2 ( .A(n9), .B(rx_ui_1_2[4]), .CI(add_263_carry[2]), .CO(
        add_263_carry[3]), .SO(rx_ui_3_8[2]) );
  FAD1X1 add_263_U1_3 ( .A(rx_ui_1_2[4]), .B(gt_647_B_3_), .CI(
        add_263_carry[3]), .CO(add_263_carry[4]), .SO(rx_ui_3_8[3]) );
  FAD1X1 add_263_U1_4 ( .A(gt_647_B_3_), .B(rx_ui_1_2[6]), .CI(
        add_263_carry[4]), .CO(add_263_carry[5]), .SO(rx_ui_3_8[4]) );
  FAD1X1 add_274_2_U1_6 ( .A(N160), .B(ui_intv_cnt[6]), .CI(add_274_2_carry[6]), .CO(add_274_2_carry[7]), .SO(N172) );
  FAD1X1 add_274_2_U1_7 ( .A(N161), .B(ui_intv_cnt[7]), .CI(add_274_2_carry[7]), .CO(add_274_2_carry[8]), .SO(N173) );
  HAD1X1 mult_274_2_U8 ( .A(symb_cnt[2]), .B(N159), .CO(mult_274_2_n7), .SO(
        N161) );
  FAD1X1 mult_274_2_U7 ( .A(symb_cnt[3]), .B(N160), .CI(mult_274_2_n7), .CO(
        mult_274_2_n6), .SO(N162) );
  FAD1X1 mult_274_2_U6 ( .A(symb_cnt[4]), .B(symb_cnt[2]), .CI(mult_274_2_n6), 
        .CO(mult_274_2_n5), .SO(N163) );
  FAD1X1 mult_274_2_U5 ( .A(symb_cnt[5]), .B(symb_cnt[3]), .CI(mult_274_2_n5), 
        .CO(mult_274_2_n4), .SO(N164) );
  FAD1X1 mult_274_2_U4 ( .A(symb_cnt[6]), .B(symb_cnt[4]), .CI(mult_274_2_n4), 
        .CO(mult_274_2_n3), .SO(N165) );
  HAD1X1 mult_274_2_U3 ( .A(mult_274_2_n3), .B(symb_cnt[5]), .CO(mult_274_2_n2), .SO(N166) );
  HAD1X1 mult_274_2_U2 ( .A(mult_274_2_n2), .B(symb_cnt[6]), .CO(N168), .SO(
        N167) );
  FAD1X1 add_274_U1_6 ( .A(N107), .B(ui_intv_cnt[6]), .CI(add_274_carry[6]), 
        .CO(add_274_carry[7]), .SO(N144) );
  FAD1X1 add_274_U1_7 ( .A(N108), .B(ui_intv_cnt[7]), .CI(add_274_carry[7]), 
        .CO(add_274_carry[8]), .SO(N145) );
  HAD1X1 mult_274_U29 ( .A(N95), .B(n296), .CO(mult_274_n7), .SO(N108) );
  FAD1X1 mult_274_U28 ( .A(N96), .B(N107), .CI(mult_274_n7), .CO(mult_274_n6), 
        .SO(N109) );
  FAD1X1 mult_274_U27 ( .A(N97), .B(N95), .CI(mult_274_n6), .CO(mult_274_n5), 
        .SO(N110) );
  FAD1X1 mult_274_U26 ( .A(N98), .B(N96), .CI(mult_274_n5), .CO(mult_274_n4), 
        .SO(N111) );
  FAD1X1 mult_274_U25 ( .A(N99), .B(N97), .CI(mult_274_n4), .CO(mult_274_n3), 
        .SO(N112) );
  FAD1X1 mult_274_U24 ( .A(N116), .B(N98), .CI(mult_274_n3), .CO(mult_274_n2), 
        .SO(N113) );
  FAD1X1 mult_274_U23 ( .A(N116), .B(N99), .CI(mult_274_n2), .CO(N115), .SO(
        N114) );
  DFFRQX1 rxtx_buf_reg_8_ ( .D(trans_buf[8]), .C(net9488), .XR(n47), .Q(
        rxtx_buf[8]) );
  DFFRQX1 rxtx_buf_reg_9_ ( .D(trans_buf[9]), .C(net9488), .XR(n47), .Q(
        rxtx_buf[9]) );
  DFFRQX1 rxtx_buf_reg_10_ ( .D(trans_buf[10]), .C(net9488), .XR(n47), .Q(
        rxtx_buf[10]) );
  DFFRQX1 rxtx_buf_reg_7_ ( .D(trans_buf[7]), .C(net9488), .XR(n47), .Q(
        rxtx_buf[7]) );
  DFFRQX1 rx_byte_pchk_reg ( .D(N356), .C(clk), .XR(n50), .Q(setsta[5]) );
  DFFRQX1 rxtx_buf_reg_1_ ( .D(trans_buf[1]), .C(net9488), .XR(n49), .Q(
        rxtx_buf[1]) );
  DFFQX1 rx_trans_8_chg_reg ( .D(n516), .C(clk), .Q(rx_trans_8_chg) );
  DFFRQX1 rxtx_buf_reg_0_ ( .D(trans_buf[0]), .C(net9488), .XR(n48), .Q(
        rxtx_buf[0]) );
  DFFRQX1 rxtx_buf_reg_2_ ( .D(trans_buf[2]), .C(net9488), .XR(n47), .Q(
        rxtx_buf[2]) );
  DFFRQX1 rxtx_buf_reg_3_ ( .D(trans_buf[3]), .C(net9488), .XR(n48), .Q(
        rxtx_buf[3]) );
  DFFRQX1 rxtx_buf_reg_5_ ( .D(trans_buf[5]), .C(net9488), .XR(n47), .Q(
        rxtx_buf[5]) );
  DFFRQX1 rxtx_buf_reg_4_ ( .D(trans_buf[4]), .C(net9488), .XR(n47), .Q(
        rxtx_buf[4]) );
  DFFRQX1 rxtx_buf_reg_6_ ( .D(trans_buf[6]), .C(net9488), .XR(n47), .Q(
        rxtx_buf[6]) );
  DFFRQX1 new_rx_sync_cnt_reg_0_ ( .D(N348), .C(clk), .XR(n41), .Q(
        new_rx_sync_cnt[0]) );
  DFFRQX1 new_rx_sync_cnt_reg_1_ ( .D(N349), .C(clk), .XR(n44), .Q(
        new_rx_sync_cnt[1]) );
  DFFSQX1 catch_sync_reg_5_ ( .D(n7), .C(net9465), .XS(n46), .Q(catch_sync[5])
         );
  DFFRQX1 us_cnt_reg_3_ ( .D(N88), .C(clk), .XR(n43), .Q(us_cnt[3]) );
  DFFRQX1 us_cnt_reg_2_ ( .D(N87), .C(clk), .XR(n45), .Q(us_cnt[2]) );
  DFFSQX1 catch_sync_reg_3_ ( .D(n14), .C(net9465), .XS(n46), .Q(catch_sync[3]) );
  DFFRQX1 catch_sync_reg_4_ ( .D(n17), .C(net9465), .XR(n48), .Q(catch_sync[4]) );
  DFFRQX1 catch_sync_reg_1_ ( .D(n13), .C(net9465), .XR(n48), .Q(catch_sync[1]) );
  DFFRQX1 catch_sync_reg_2_ ( .D(ui_intv_cnt[2]), .C(net9465), .XR(n48), .Q(
        catch_sync[2]) );
  DFFRQX1 us_cnt_reg_1_ ( .D(n461), .C(clk), .XR(srstz), .Q(us_cnt[1]) );
  DFFRQX1 us_cnt_reg_0_ ( .D(N85), .C(clk), .XR(n47), .Q(us_cnt[0]) );
  DFFRQX1 sync_length_reg_1_ ( .D(N261), .C(net9483), .XR(n49), .Q(N363) );
  DFFRQX1 sync_length_reg_0_ ( .D(N260), .C(net9483), .XR(n49), .Q(N362) );
  DFFRQX1 catch_sync_reg_0_ ( .D(ui_intv_cnt[0]), .C(net9465), .XR(n48), .Q(
        catch_sync[0]) );
  DFFRQX1 ui_intv_cnt_reg_0_ ( .D(net9480), .C(net9483), .XR(n48), .Q(
        ui_intv_cnt[0]) );
  DFFRQX1 symb_cnt_reg_4_ ( .D(N1014), .C(net9498), .XR(n50), .Q(symb_cnt[4])
         );
  DFFRQX1 ui_intv_cnt_reg_1_ ( .D(net9477), .C(net9483), .XR(n48), .Q(
        ui_intv_cnt[1]) );
  DFFRQX1 symb_cnt_reg_6_ ( .D(N1016), .C(net9498), .XR(n49), .Q(symb_cnt[6])
         );
  DFFRQX1 symb_cnt_reg_5_ ( .D(N1015), .C(net9498), .XR(n50), .Q(symb_cnt[5])
         );
  DFFRQX1 ui_intv_cnt_reg_6_ ( .D(net9472), .C(net9483), .XR(n49), .Q(
        ui_intv_cnt[6]) );
  DFFRQX1 ui_intv_cnt_reg_7_ ( .D(net9469), .C(net9483), .XR(n49), .Q(
        ui_intv_cnt[7]) );
  DFFRQX1 ui_intv_cnt_reg_2_ ( .D(net9476), .C(net9483), .XR(n48), .Q(
        ui_intv_cnt[2]) );
  DFFRQX1 ui_intv_cnt_reg_5_ ( .D(net9473), .C(net9483), .XR(n49), .Q(
        ui_intv_cnt[5]) );
  DFFRQX1 ui_intv_cnt_reg_3_ ( .D(net9475), .C(net9483), .XR(n48), .Q(N141) );
  DFFRQX1 ui_intv_cnt_reg_4_ ( .D(net9474), .C(net9483), .XR(n49), .Q(N142) );
  DFFRQX1 symb_cnt_reg_3_ ( .D(N1013), .C(net9498), .XR(n50), .Q(symb_cnt[3])
         );
  DFFRQX1 symb_cnt_reg_2_ ( .D(N1012), .C(net9498), .XR(n50), .Q(symb_cnt[2])
         );
  DFFRQX1 symb_cnt_reg_1_ ( .D(N1011), .C(net9498), .XR(n50), .Q(N160) );
  DFFRQX1 symb_cnt_reg_0_ ( .D(N1010), .C(net9498), .XR(n50), .Q(N159) );
  DFFRQX1 rxtx_buf_reg_11_ ( .D(trans_buf[11]), .C(net9488), .XR(n49), .Q(
        tx_dat) );
  DFFSQX1 tx_dbuf_keep_empty_reg ( .D(N444), .C(clk), .XS(n47), .Q(r_ctl[7])
         );
  DFFRQX1 fcp_state_reg_2_ ( .D(N1008), .C(net9493), .XR(n50), .Q(fcp_state[2]) );
  DFFRQX1 fcp_state_reg_1_ ( .D(N1007), .C(net9493), .XR(n50), .Q(fcp_state[1]) );
  DFFRQX1 fcp_state_reg_0_ ( .D(N1006), .C(net9493), .XR(n50), .Q(fcp_state[0]) );
  DFFRQX1 fcp_state_reg_3_ ( .D(N1009), .C(net9493), .XR(n49), .Q(fcp_state[3]) );
  NOR2X1 U3 ( .A(sub_423_carry_5_), .B(rx_ui_1_2[6]), .Y(n1) );
  INVX1 U4 ( .A(n276), .Y(n2) );
  INVX1 U5 ( .A(n188), .Y(n3) );
  INVX1 U6 ( .A(n297), .Y(n4) );
  INVX1 U7 ( .A(r_ctl[0]), .Y(n5) );
  INVX1 U8 ( .A(n360), .Y(n6) );
  BUFX3 U9 ( .A(ui_intv_cnt[5]), .Y(n7) );
  INVX1 U10 ( .A(n137), .Y(n8) );
  MUX2IX1 U11 ( .D0(catch_sync[2]), .D1(r_tui[4]), .S(n92), .Y(N326) );
  INVX1 U12 ( .A(N326), .Y(n9) );
  INVX1 U13 ( .A(N326), .Y(n10) );
  INVX1 U14 ( .A(n333), .Y(n11) );
  INVX1 U15 ( .A(n186), .Y(n22) );
  INVX1 U16 ( .A(n22), .Y(n12) );
  INVX1 U17 ( .A(n86), .Y(n13) );
  INVX1 U18 ( .A(n66), .Y(n14) );
  BUFX3 U19 ( .A(n152), .Y(n15) );
  INVX1 U20 ( .A(n364), .Y(n16) );
  INVX1 U21 ( .A(n187), .Y(n17) );
  INVX1 U22 ( .A(n296), .Y(n18) );
  INVX1 U23 ( .A(n51), .Y(n46) );
  INVX1 U24 ( .A(n51), .Y(n47) );
  INVX1 U25 ( .A(n51), .Y(n48) );
  INVX1 U26 ( .A(n51), .Y(n49) );
  INVX1 U27 ( .A(n51), .Y(n50) );
  INVX1 U28 ( .A(n51), .Y(n45) );
  INVX1 U29 ( .A(n51), .Y(n43) );
  INVX1 U30 ( .A(n51), .Y(n44) );
  INVX1 U31 ( .A(n51), .Y(n41) );
  INVX1 U32 ( .A(srstz), .Y(n51) );
  INVX1 U33 ( .A(n40), .Y(n39) );
  INVX1 U34 ( .A(n33), .Y(n25) );
  INVX1 U35 ( .A(n38), .Y(n37) );
  INVX1 U36 ( .A(r_wdat[2]), .Y(n33) );
  INVX1 U37 ( .A(r_wdat[7]), .Y(n40) );
  INVX1 U38 ( .A(r_wdat[6]), .Y(n38) );
  INVX1 U39 ( .A(r_wdat[5]), .Y(n36) );
  INVX1 U40 ( .A(r_wdat[4]), .Y(n35) );
  INVX1 U41 ( .A(r_wdat[3]), .Y(n34) );
  INVX1 U42 ( .A(r_wdat[0]), .Y(n23) );
  INVX1 U43 ( .A(r_wdat[1]), .Y(n24) );
  NAND21X1 U44 ( .B(ui_by_ping[5]), .A(n93), .Y(n97) );
  INVX1 U45 ( .A(n134), .Y(n123) );
  XOR2X1 U46 ( .A(sub_423_carry_5_), .B(rx_ui_1_2[6]), .Y(n19) );
  NOR2X1 U47 ( .A(n152), .B(n151), .Y(n122) );
  INVX1 U48 ( .A(n364), .Y(N325) );
  GEN2XL U49 ( .D(n88), .E(n187), .C(n87), .B(n188), .A(n189), .Y(n186) );
  INVX1 U50 ( .A(n277), .Y(gt_647_B_3_) );
  INVX1 U51 ( .A(n276), .Y(n80) );
  INVX1 U52 ( .A(n361), .Y(rx_ui_1_2[4]) );
  INVX1 U53 ( .A(n61), .Y(n68) );
  INVX1 U54 ( .A(n360), .Y(rx_ui_1_2[6]) );
  NAND2X1 U55 ( .A(n259), .B(n333), .Y(n246) );
  INVX1 U56 ( .A(ui_intv_cnt[5]), .Y(n88) );
  NOR3XL U57 ( .A(n164), .B(r_ctl[7]), .C(n165), .Y(n152) );
  INVX1 U58 ( .A(n58), .Y(n67) );
  NAND4X1 U59 ( .A(n446), .B(n447), .C(n448), .D(n449), .Y(n165) );
  INVX1 U60 ( .A(r_tui[5]), .Y(adp_tx_ui_5_) );
  INVX1 U61 ( .A(symb_cnt[2]), .Y(n308) );
  INVX1 U62 ( .A(N141), .Y(n66) );
  INVX1 U63 ( .A(r_ctl[0]), .Y(n121) );
  BUFX3 U64 ( .A(r_ctl[6]), .Y(tx_en) );
  BUFX3 U65 ( .A(ff_idn), .Y(r_ctl[5]) );
  AND2X1 U66 ( .A(catch_ping[15]), .B(add_277_carry[11]), .Y(ui_by_ping[12])
         );
  XOR2X1 U67 ( .A(add_277_carry[11]), .B(catch_ping[15]), .Y(ui_by_ping[11])
         );
  AND2X1 U68 ( .A(add_277_carry[10]), .B(catch_ping[14]), .Y(add_277_carry[11]) );
  XOR2X1 U69 ( .A(add_277_carry[10]), .B(catch_ping[14]), .Y(ui_by_ping[10])
         );
  AND2X1 U70 ( .A(add_277_carry[9]), .B(catch_ping[13]), .Y(add_277_carry[10])
         );
  XOR2X1 U71 ( .A(add_277_carry[9]), .B(catch_ping[13]), .Y(ui_by_ping[9]) );
  AND2X1 U72 ( .A(add_277_carry[8]), .B(catch_ping[12]), .Y(add_277_carry[9])
         );
  XOR2X1 U74 ( .A(add_277_carry[8]), .B(catch_ping[12]), .Y(ui_by_ping[8]) );
  AND2X1 U75 ( .A(add_277_carry[7]), .B(catch_ping[11]), .Y(add_277_carry[8])
         );
  XOR2X1 U76 ( .A(add_277_carry[7]), .B(catch_ping[11]), .Y(ui_by_ping[7]) );
  AND2X1 U77 ( .A(N168), .B(add_274_2_carry[14]), .Y(N181) );
  XOR2X1 U78 ( .A(add_274_2_carry[14]), .B(N168), .Y(N180) );
  AND2X1 U79 ( .A(N167), .B(add_274_2_carry[13]), .Y(add_274_2_carry[14]) );
  XOR2X1 U80 ( .A(add_274_2_carry[13]), .B(N167), .Y(N179) );
  AND2X1 U81 ( .A(N166), .B(add_274_2_carry[12]), .Y(add_274_2_carry[13]) );
  XOR2X1 U82 ( .A(add_274_2_carry[12]), .B(N166), .Y(N178) );
  AND2X1 U83 ( .A(N165), .B(add_274_2_carry[11]), .Y(add_274_2_carry[12]) );
  XOR2X1 U84 ( .A(add_274_2_carry[11]), .B(N165), .Y(N177) );
  XOR2X1 U85 ( .A(N116), .B(add_274_carry[15]), .Y(N153) );
  AND2X1 U86 ( .A(N115), .B(add_274_carry[14]), .Y(add_274_carry[15]) );
  XOR2X1 U87 ( .A(add_274_carry[14]), .B(N115), .Y(N152) );
  AND2X1 U88 ( .A(N114), .B(add_274_carry[13]), .Y(add_274_carry[14]) );
  XOR2X1 U89 ( .A(add_274_carry[13]), .B(N114), .Y(N151) );
  AND2X1 U90 ( .A(N113), .B(add_274_carry[12]), .Y(add_274_carry[13]) );
  XOR2X1 U91 ( .A(add_274_carry[12]), .B(N113), .Y(N150) );
  AND2X1 U92 ( .A(N112), .B(add_274_carry[11]), .Y(add_274_carry[12]) );
  XOR2X1 U93 ( .A(add_274_carry[11]), .B(N112), .Y(N149) );
  XNOR2XL U94 ( .A(ui_by_ping[6]), .B(ui_by_ping[5]), .Y(N192) );
  AND2X1 U95 ( .A(add_277_carry[6]), .B(catch_ping[10]), .Y(add_277_carry[7])
         );
  XOR2X1 U96 ( .A(add_277_carry[6]), .B(catch_ping[10]), .Y(ui_by_ping[6]) );
  AND2X1 U97 ( .A(add_277_carry[5]), .B(catch_ping[9]), .Y(add_277_carry[6])
         );
  XOR2X1 U98 ( .A(add_277_carry[5]), .B(catch_ping[9]), .Y(ui_by_ping[5]) );
  AND2X1 U99 ( .A(catch_ping[8]), .B(add_277_carry[4]), .Y(add_277_carry[5])
         );
  XOR2X1 U100 ( .A(add_277_carry[4]), .B(catch_ping[8]), .Y(N190) );
  AND2X1 U101 ( .A(catch_ping[7]), .B(add_277_carry[3]), .Y(add_277_carry[4])
         );
  XOR2X1 U102 ( .A(add_277_carry[3]), .B(catch_ping[7]), .Y(N189) );
  AND2X1 U103 ( .A(catch_ping[6]), .B(add_277_carry[2]), .Y(add_277_carry[3])
         );
  XOR2X1 U104 ( .A(add_277_carry[2]), .B(catch_ping[6]), .Y(N188) );
  AND2X1 U105 ( .A(catch_ping[5]), .B(add_277_carry[1]), .Y(add_277_carry[2])
         );
  XOR2X1 U106 ( .A(add_277_carry[1]), .B(catch_ping[5]), .Y(N187) );
  AND2X1 U107 ( .A(catch_ping[3]), .B(catch_ping[4]), .Y(add_277_carry[1]) );
  XOR2X1 U108 ( .A(catch_ping[4]), .B(catch_ping[3]), .Y(N186) );
  AND2X1 U109 ( .A(N164), .B(add_274_2_carry[10]), .Y(add_274_2_carry[11]) );
  XOR2X1 U110 ( .A(add_274_2_carry[10]), .B(N164), .Y(N176) );
  AND2X1 U111 ( .A(N163), .B(add_274_2_carry[9]), .Y(add_274_2_carry[10]) );
  XOR2X1 U112 ( .A(add_274_2_carry[9]), .B(N163), .Y(N175) );
  AND2X1 U113 ( .A(N162), .B(add_274_2_carry[8]), .Y(add_274_2_carry[9]) );
  XOR2X1 U114 ( .A(add_274_2_carry[8]), .B(N162), .Y(N174) );
  AND2X1 U115 ( .A(ui_intv_cnt[5]), .B(N159), .Y(add_274_2_carry[6]) );
  XOR2X1 U116 ( .A(N159), .B(ui_intv_cnt[5]), .Y(N171) );
  AND2X1 U117 ( .A(N111), .B(add_274_carry[10]), .Y(add_274_carry[11]) );
  XOR2X1 U118 ( .A(add_274_carry[10]), .B(N111), .Y(N148) );
  AND2X1 U119 ( .A(N110), .B(add_274_carry[9]), .Y(add_274_carry[10]) );
  XOR2X1 U120 ( .A(add_274_carry[9]), .B(N110), .Y(N147) );
  AND2X1 U121 ( .A(N109), .B(add_274_carry[8]), .Y(add_274_carry[9]) );
  XOR2X1 U122 ( .A(add_274_carry[8]), .B(N109), .Y(N146) );
  AND2X1 U123 ( .A(ui_intv_cnt[5]), .B(n296), .Y(add_274_carry[6]) );
  XOR2X1 U124 ( .A(n296), .B(ui_intv_cnt[5]), .Y(N143) );
  AND2X1 U125 ( .A(n6), .B(add_264_carry[6]), .Y(rx_ui_5_8[7]) );
  XOR2X1 U126 ( .A(add_264_carry[6]), .B(n6), .Y(rx_ui_5_8[6]) );
  AND2X1 U127 ( .A(add_264_carry[5]), .B(gt_647_B_3_), .Y(add_264_carry[6]) );
  XOR2X1 U128 ( .A(add_264_carry[5]), .B(gt_647_B_3_), .Y(rx_ui_5_8[5]) );
  AND2X1 U129 ( .A(add_264_A_0_), .B(N325), .Y(add_264_carry[1]) );
  XOR2X1 U130 ( .A(add_264_A_0_), .B(n16), .Y(rx_ui_5_8[0]) );
  OR2X1 U131 ( .A(rx_ui_1_2[4]), .B(gt_647_B_3_), .Y(sub_423_carry_5_) );
  XNOR2XL U132 ( .A(rx_ui_1_2[4]), .B(gt_647_B_3_), .Y(N328) );
  AND2X1 U133 ( .A(rx_ui_1_2[6]), .B(add_423_carry_5_), .Y(N338) );
  XOR2X1 U134 ( .A(add_423_carry_5_), .B(rx_ui_1_2[6]), .Y(N337) );
  AND2X1 U135 ( .A(gt_647_B_3_), .B(rx_ui_1_2[4]), .Y(add_423_carry_5_) );
  XOR2X1 U136 ( .A(n231), .B(gt_647_B_3_), .Y(N336) );
  AND2X1 U137 ( .A(rx_ui_1_2[6]), .B(add_263_carry[5]), .Y(rx_ui_3_8[6]) );
  XOR2X1 U138 ( .A(add_263_carry[5]), .B(rx_ui_1_2[6]), .Y(rx_ui_3_8[5]) );
  AND2X1 U139 ( .A(N324), .B(N325), .Y(add_263_carry[1]) );
  XOR2X1 U140 ( .A(N324), .B(N325), .Y(rx_ui_3_8[0]) );
  AND2X1 U141 ( .A(N363), .B(N362), .Y(N419) );
  XOR2X1 U142 ( .A(N362), .B(N363), .Y(N418) );
  XNOR2XL U143 ( .A(r_tui[6]), .B(add_282_carry_7_), .Y(adp_tx_ui_7_) );
  AND2X1 U144 ( .A(r_tui[5]), .B(r_tui[6]), .Y(add_282_carry_7_) );
  XOR2X1 U145 ( .A(r_tui[5]), .B(r_tui[6]), .Y(adp_tx_ui_6_) );
  AND2X1 U146 ( .A(ui_intv_cnt[0]), .B(N219), .Y(N1252) );
  AND2X1 U147 ( .A(n13), .B(N219), .Y(N1253) );
  AND2X1 U148 ( .A(ui_intv_cnt[2]), .B(N219), .Y(N1254) );
  AND2X1 U149 ( .A(n14), .B(N219), .Y(N1255) );
  AND2X1 U150 ( .A(n17), .B(N219), .Y(N1256) );
  AND2X1 U151 ( .A(n7), .B(N219), .Y(N1257) );
  AND2X1 U152 ( .A(ui_intv_cnt[6]), .B(N219), .Y(N1258) );
  AND2X1 U153 ( .A(N219), .B(ui_intv_cnt[7]), .Y(N1259) );
  OR2X1 U154 ( .A(N160), .B(N159), .Y(n52) );
  OAI21BBX1 U155 ( .A(N159), .B(N160), .C(n52), .Y(N107) );
  OR2X1 U156 ( .A(n52), .B(symb_cnt[2]), .Y(n53) );
  OAI21BBX1 U157 ( .A(n52), .B(symb_cnt[2]), .C(n53), .Y(N95) );
  OR2X1 U158 ( .A(n53), .B(symb_cnt[3]), .Y(n54) );
  OAI21BBX1 U159 ( .A(n53), .B(symb_cnt[3]), .C(n54), .Y(N96) );
  OR2X1 U160 ( .A(n54), .B(symb_cnt[4]), .Y(n55) );
  OAI21BBX1 U161 ( .A(n54), .B(symb_cnt[4]), .C(n55), .Y(N97) );
  XNOR2XL U162 ( .A(n55), .B(symb_cnt[5]), .Y(N98) );
  OR2X1 U163 ( .A(symb_cnt[5]), .B(n55), .Y(n56) );
  NOR3XL U164 ( .A(symb_cnt[5]), .B(symb_cnt[6]), .C(n55), .Y(N116) );
  AO21X1 U165 ( .B(n56), .C(symb_cnt[6]), .A(N116), .Y(N99) );
  NOR2X1 U166 ( .A(n19), .B(ui_intv_cnt[5]), .Y(n61) );
  AOI32X1 U167 ( .A(n68), .B(N336), .C(N142), .D(ui_intv_cnt[5]), .E(n19), .Y(
        n65) );
  AND2X1 U168 ( .A(n361), .B(n66), .Y(n60) );
  OAI32X1 U169 ( .A(n233), .B(n10), .C(n60), .D(n361), .E(n66), .Y(n58) );
  AOI22BXL U170 ( .B(ui_intv_cnt[1]), .A(N325), .D(ui_intv_cnt[0]), .C(N324), 
        .Y(n57) );
  AOI211X1 U171 ( .C(ui_intv_cnt[1]), .D(n364), .A(n58), .B(n57), .Y(n59) );
  GEN2XL U172 ( .D(n10), .E(n233), .C(n60), .B(n67), .A(n59), .Y(n62) );
  AOI211X1 U173 ( .C(N328), .D(n187), .A(n62), .B(n61), .Y(n63) );
  NOR3XL U174 ( .A(n63), .B(ui_intv_cnt[7]), .C(ui_intv_cnt[6]), .Y(n64) );
  AOI21X1 U175 ( .B(n65), .C(n64), .A(n1), .Y(N331) );
  OAI21X1 U176 ( .B(n69), .C(n70), .A(n71), .Y(upd_dbuf_en) );
  NAND4X1 U177 ( .A(n72), .B(n73), .C(n74), .D(n75), .Y(n70) );
  XNOR2XL U178 ( .A(ui_intv_cnt[2]), .B(rx_ui_5_8[2]), .Y(n75) );
  NOR2X1 U179 ( .A(n76), .B(n77), .Y(n74) );
  XNOR2XL U180 ( .A(rx_ui_5_8[0]), .B(n78), .Y(n77) );
  XNOR2XL U181 ( .A(rx_ui_5_8[3]), .B(n66), .Y(n76) );
  XNOR2XL U182 ( .A(n17), .B(rx_ui_5_8[4]), .Y(n73) );
  XNOR2XL U183 ( .A(ui_intv_cnt[7]), .B(rx_ui_5_8[7]), .Y(n72) );
  NAND4X1 U184 ( .A(n79), .B(n80), .C(n81), .D(n82), .Y(n69) );
  NOR3XL U185 ( .A(n83), .B(n84), .C(n85), .Y(n82) );
  XNOR2XL U186 ( .A(rx_ui_5_8[1]), .B(n86), .Y(n85) );
  XNOR2XL U187 ( .A(rx_ui_5_8[6]), .B(n87), .Y(n84) );
  XNOR2XL U188 ( .A(rx_ui_5_8[5]), .B(n88), .Y(n83) );
  MUX2X1 U189 ( .D0(n39), .D1(rxtx_buf[7]), .S(n71), .Y(upd_dbuf[7]) );
  MUX2X1 U190 ( .D0(n37), .D1(rxtx_buf[6]), .S(n71), .Y(upd_dbuf[6]) );
  MUX2X1 U191 ( .D0(r_wdat[5]), .D1(rxtx_buf[5]), .S(n71), .Y(upd_dbuf[5]) );
  MUX2X1 U192 ( .D0(r_wdat[4]), .D1(rxtx_buf[4]), .S(n71), .Y(upd_dbuf[4]) );
  MUX2X1 U193 ( .D0(r_wdat[3]), .D1(rxtx_buf[3]), .S(n71), .Y(upd_dbuf[3]) );
  INVX1 U194 ( .A(r_wr[3]), .Y(n71) );
  MUX2IX1 U195 ( .D0(n89), .D1(n33), .S(r_wr[3]), .Y(upd_dbuf[2]) );
  MUX2IX1 U196 ( .D0(n90), .D1(n24), .S(r_wr[3]), .Y(upd_dbuf[1]) );
  MUX2IX1 U197 ( .D0(n91), .D1(n23), .S(r_wr[3]), .Y(upd_dbuf[0]) );
  MUX2IX1 U198 ( .D0(n92), .D1(n40), .S(r_wr[4]), .Y(tui_wdat[7]) );
  OAI21BBX1 U199 ( .A(N192), .B(n93), .C(n94), .Y(tui_wdat[6]) );
  MUX2IX1 U200 ( .D0(n95), .D1(n37), .S(r_wr[4]), .Y(n94) );
  OAI211X1 U201 ( .C(n36), .D(n96), .A(n97), .B(n98), .Y(tui_wdat[5]) );
  OAI211X1 U202 ( .C(n35), .D(n96), .A(n99), .B(n98), .Y(tui_wdat[4]) );
  NAND2X1 U203 ( .A(N190), .B(n93), .Y(n99) );
  OAI211X1 U204 ( .C(n34), .D(n96), .A(n100), .B(n98), .Y(tui_wdat[3]) );
  NAND2X1 U205 ( .A(N189), .B(n93), .Y(n100) );
  OAI2B11X1 U206 ( .D(n93), .C(n101), .A(n98), .B(n102), .Y(tui_wdat[2]) );
  MUX2IX1 U207 ( .D0(n95), .D1(n25), .S(r_wr[4]), .Y(n102) );
  NAND2X1 U208 ( .A(n103), .B(n96), .Y(n98) );
  INVX1 U209 ( .A(N188), .Y(n101) );
  ENOX1 U210 ( .A(n24), .B(n96), .C(N187), .D(n93), .Y(tui_wdat[1]) );
  ENOX1 U211 ( .A(n23), .B(n96), .C(N186), .D(n93), .Y(tui_wdat[0]) );
  NOR3XL U212 ( .A(n95), .B(r_wr[4]), .C(n103), .Y(n93) );
  NAND43X1 U213 ( .B(ui_by_ping[8]), .C(ui_by_ping[9]), .D(ui_by_ping[12]), 
        .A(n104), .Y(n103) );
  AOI211X1 U214 ( .C(n105), .D(n106), .A(ui_by_ping[11]), .B(ui_by_ping[10]), 
        .Y(n104) );
  OAI21BX1 U215 ( .C(N190), .B(n107), .A(n108), .Y(n106) );
  OAI21BX1 U216 ( .C(N189), .B(n109), .A(n108), .Y(n105) );
  NAND21X1 U217 ( .B(n107), .A(ui_by_ping[5]), .Y(n108) );
  NAND2X1 U218 ( .A(ui_by_ping[7]), .B(ui_by_ping[6]), .Y(n107) );
  OAI21X1 U219 ( .B(N186), .C(N187), .A(N188), .Y(n109) );
  AND2X1 U220 ( .A(n110), .B(n111), .Y(n95) );
  NOR4XL U221 ( .A(ui_by_ping[9]), .B(ui_by_ping[8]), .C(ui_by_ping[7]), .D(
        ui_by_ping[12]), .Y(n111) );
  AOI211X1 U222 ( .C(n112), .D(ui_by_ping[6]), .A(ui_by_ping[11]), .B(
        ui_by_ping[10]), .Y(n110) );
  INVX1 U223 ( .A(n113), .Y(n112) );
  OAI31XL U224 ( .A(N189), .B(N190), .C(N188), .D(ui_by_ping[5]), .Y(n113) );
  OAI31XL U225 ( .A(n114), .B(n115), .C(n116), .D(n96), .Y(tui_upd) );
  INVX1 U226 ( .A(r_wr[4]), .Y(n96) );
  INVX1 U227 ( .A(n117), .Y(n116) );
  NAND2X1 U228 ( .A(n118), .B(n119), .Y(trans_buf[9]) );
  AOI22X1 U229 ( .A(n120), .B(n121), .C(rxtx_buf[8]), .D(n122), .Y(n118) );
  AO2222XL U230 ( .A(n122), .B(rxtx_buf[7]), .C(n123), .D(n124), .E(n125), .F(
        n121), .G(n126), .H(n127), .Y(trans_buf[8]) );
  AO2222XL U231 ( .A(n122), .B(rxtx_buf[6]), .C(n123), .D(n127), .E(n128), .F(
        n121), .G(n129), .H(n120), .Y(trans_buf[7]) );
  AO2222XL U232 ( .A(n122), .B(rxtx_buf[5]), .C(n123), .D(n120), .E(n130), .F(
        n121), .G(n129), .H(n125), .Y(trans_buf[6]) );
  AO2222XL U233 ( .A(n122), .B(rxtx_buf[4]), .C(n131), .D(n121), .E(n123), .F(
        n125), .G(n129), .H(n128), .Y(trans_buf[5]) );
  AO2222XL U234 ( .A(n8), .B(rxtx_buf[3]), .C(n132), .D(n121), .E(n123), .F(
        n128), .G(n129), .H(n130), .Y(trans_buf[4]) );
  OAI222XL U235 ( .A(n133), .B(n134), .C(n135), .D(n136), .E(n89), .F(n137), 
        .Y(trans_buf[3]) );
  INVX1 U236 ( .A(rxtx_buf[2]), .Y(n89) );
  OAI222XL U237 ( .A(n135), .B(n134), .C(n138), .D(n136), .E(n90), .F(n137), 
        .Y(trans_buf[2]) );
  INVX1 U238 ( .A(rxtx_buf[1]), .Y(n90) );
  OAI21X1 U239 ( .B(n91), .C(n137), .A(n139), .Y(trans_buf[1]) );
  AOI32X1 U240 ( .A(n126), .B(n140), .C(n141), .D(n123), .E(n132), .Y(n139) );
  INVX1 U241 ( .A(rxtx_buf[0]), .Y(n91) );
  NAND2X1 U242 ( .A(n142), .B(n119), .Y(trans_buf[11]) );
  MUX2IX1 U243 ( .D0(n129), .D1(n123), .S(n143), .Y(n119) );
  AOI22X1 U244 ( .A(n124), .B(n121), .C(rxtx_buf[10]), .D(n122), .Y(n142) );
  NAND2X1 U245 ( .A(n144), .B(n145), .Y(trans_buf[10]) );
  MUX2IX1 U246 ( .D0(n123), .D1(n126), .S(n143), .Y(n145) );
  INVX1 U247 ( .A(n136), .Y(n126) );
  NAND2X1 U248 ( .A(n129), .B(n137), .Y(n136) );
  NOR2X1 U249 ( .A(n121), .B(n123), .Y(n129) );
  AOI22X1 U250 ( .A(n127), .B(n121), .C(rxtx_buf[9]), .D(n122), .Y(n144) );
  AO33X1 U251 ( .A(r_ctl[5]), .B(n146), .C(n122), .D(n141), .E(n140), .F(n123), 
        .Y(trans_buf[0]) );
  XNOR2XL U252 ( .A(n147), .B(n148), .Y(n141) );
  XNOR2XL U253 ( .A(n149), .B(n150), .Y(n148) );
  XNOR2XL U254 ( .A(n130), .B(n124), .Y(n150) );
  INVX1 U255 ( .A(n143), .Y(n124) );
  AOI22X1 U256 ( .A(n39), .B(n151), .C(n152), .D(r_dat[7]), .Y(n143) );
  INVX1 U257 ( .A(n133), .Y(n130) );
  AOI22X1 U258 ( .A(n25), .B(n151), .C(r_dat[2]), .D(n152), .Y(n133) );
  XNOR2XL U259 ( .A(n131), .B(n132), .Y(n149) );
  INVX1 U260 ( .A(n138), .Y(n132) );
  AOI22X1 U261 ( .A(r_wdat[0]), .B(n151), .C(r_dat[0]), .D(n152), .Y(n138) );
  INVX1 U262 ( .A(n135), .Y(n131) );
  AOI22X1 U263 ( .A(r_wdat[1]), .B(n151), .C(r_dat[1]), .D(n152), .Y(n135) );
  XNOR2XL U264 ( .A(n153), .B(n154), .Y(n147) );
  XNOR2XL U265 ( .A(n127), .B(n120), .Y(n154) );
  ENOX1 U266 ( .A(n36), .B(n155), .C(r_dat[5]), .D(n152), .Y(n120) );
  ENOX1 U267 ( .A(n38), .B(n155), .C(r_dat[6]), .D(n152), .Y(n127) );
  XNOR2XL U268 ( .A(n128), .B(n125), .Y(n153) );
  ENOX1 U269 ( .A(n35), .B(n155), .C(r_dat[4]), .D(n152), .Y(n125) );
  ENOX1 U270 ( .A(n34), .B(n155), .C(r_dat[3]), .D(n152), .Y(n128) );
  NOR3XL U271 ( .A(n156), .B(n157), .C(n158), .Y(setsta[6]) );
  NAND3X1 U272 ( .A(ff_chg), .B(n159), .C(ff_idn), .Y(n156) );
  INVX1 U273 ( .A(n160), .Y(setsta[4]) );
  NOR32XL U274 ( .B(new_rx_sync_cnt[1]), .C(n161), .A(n162), .Y(setsta[3]) );
  NOR3XL U275 ( .A(n163), .B(n164), .C(n165), .Y(setsta[0]) );
  AOI21BBXL U276 ( .B(us_cnt[1]), .C(us_cnt[0]), .A(n166), .Y(n461) );
  OAI2B11X1 U277 ( .D(N221), .C(n167), .A(n168), .B(n169), .Y(net9480) );
  AND2X1 U278 ( .A(N222), .B(n170), .Y(net9477) );
  AND2X1 U279 ( .A(N223), .B(n170), .Y(net9476) );
  AND2X1 U280 ( .A(N224), .B(n170), .Y(net9475) );
  ENOX1 U281 ( .A(n171), .B(n168), .C(N225), .D(n170), .Y(net9474) );
  AND2X1 U282 ( .A(N226), .B(n170), .Y(net9473) );
  ENOX1 U283 ( .A(n171), .B(n168), .C(N227), .D(n170), .Y(net9472) );
  AND2X1 U284 ( .A(N228), .B(n170), .Y(net9469) );
  AND3X1 U285 ( .A(n81), .B(n168), .C(n169), .Y(n170) );
  INVX1 U286 ( .A(n172), .Y(N324) );
  NOR4XL U287 ( .A(n173), .B(n174), .C(n114), .D(n175), .Y(n525) );
  NAND21X1 U288 ( .B(n176), .A(n177), .Y(n174) );
  INVX1 U289 ( .A(n178), .Y(n517) );
  MUX2IX1 U290 ( .D0(n179), .D1(ff_chg), .S(rx_trans_8_chg), .Y(n516) );
  NAND2X1 U291 ( .A(n180), .B(n79), .Y(n179) );
  NAND4X1 U292 ( .A(n181), .B(n182), .C(n183), .D(n184), .Y(intr) );
  AOI22X1 U293 ( .A(r_msk[0]), .B(r_irq[0]), .C(r_msk[1]), .D(r_irq[1]), .Y(
        n184) );
  AOI22X1 U294 ( .A(r_msk[2]), .B(r_irq[2]), .C(r_msk[3]), .D(r_irq[3]), .Y(
        n183) );
  AOI22X1 U295 ( .A(r_msk[4]), .B(r_irq[4]), .C(r_msk[5]), .D(r_irq[5]), .Y(
        n182) );
  AOI22X1 U296 ( .A(r_msk[6]), .B(r_irq[6]), .C(r_msk[7]), .D(r_irq[7]), .Y(
        n181) );
  NOR2X1 U297 ( .A(n40), .B(n185), .Y(clrsta[7]) );
  NOR2X1 U298 ( .A(n38), .B(n185), .Y(clrsta[6]) );
  NOR2X1 U299 ( .A(n36), .B(n185), .Y(clrsta[5]) );
  NOR2X1 U300 ( .A(n35), .B(n185), .Y(clrsta[4]) );
  NOR2X1 U301 ( .A(n34), .B(n185), .Y(clrsta[3]) );
  NOR2X1 U302 ( .A(n33), .B(n185), .Y(clrsta[2]) );
  NOR2X1 U303 ( .A(n24), .B(n185), .Y(clrsta[1]) );
  NOR2X1 U304 ( .A(n23), .B(n185), .Y(clrsta[0]) );
  INVX1 U305 ( .A(r_wr[1]), .Y(n185) );
  MUX2X1 U306 ( .D0(N147), .D1(N175), .S(n12), .Y(catch_ping[9]) );
  MUX2X1 U307 ( .D0(N146), .D1(N174), .S(n12), .Y(catch_ping[8]) );
  MUX2X1 U308 ( .D0(N145), .D1(N173), .S(n12), .Y(catch_ping[7]) );
  MUX2X1 U309 ( .D0(N144), .D1(N172), .S(n12), .Y(catch_ping[6]) );
  MUX2X1 U310 ( .D0(N143), .D1(N171), .S(n186), .Y(catch_ping[5]) );
  MUX2X1 U311 ( .D0(N142), .D1(N142), .S(n186), .Y(catch_ping[4]) );
  MUX2X1 U312 ( .D0(N141), .D1(N141), .S(n186), .Y(catch_ping[3]) );
  MUX2X1 U313 ( .D0(N153), .D1(N181), .S(n12), .Y(catch_ping[15]) );
  MUX2X1 U314 ( .D0(N152), .D1(N180), .S(n12), .Y(catch_ping[14]) );
  MUX2X1 U315 ( .D0(N151), .D1(N179), .S(n12), .Y(catch_ping[13]) );
  MUX2X1 U316 ( .D0(N150), .D1(N178), .S(n12), .Y(catch_ping[12]) );
  MUX2X1 U317 ( .D0(N149), .D1(N177), .S(n12), .Y(catch_ping[11]) );
  MUX2X1 U318 ( .D0(N148), .D1(N176), .S(n12), .Y(catch_ping[10]) );
  MUX2IX1 U319 ( .D0(n190), .D1(n166), .S(us_cnt[3]), .Y(N88) );
  NAND3X1 U320 ( .A(n191), .B(n192), .C(us_cnt[2]), .Y(n190) );
  MUX2IX1 U321 ( .D0(n193), .D1(n166), .S(us_cnt[2]), .Y(N87) );
  NAND2X1 U322 ( .A(n191), .B(n194), .Y(n166) );
  NAND2X1 U323 ( .A(n191), .B(n192), .Y(n193) );
  NOR21XL U324 ( .B(n191), .A(us_cnt[0]), .Y(N85) );
  NOR2X1 U325 ( .A(n195), .B(n81), .Y(n191) );
  AOI21X1 U326 ( .B(n163), .C(n178), .A(r_wr[3]), .Y(N444) );
  OAI211X1 U327 ( .C(n196), .D(n197), .A(n198), .B(n199), .Y(n178) );
  AOI211X1 U328 ( .C(n200), .D(n201), .A(n18), .B(n146), .Y(n199) );
  INVX1 U329 ( .A(n202), .Y(n200) );
  NOR2X1 U330 ( .A(n160), .B(n203), .Y(N356) );
  XNOR2XL U331 ( .A(rxtx_buf[7]), .B(n204), .Y(n203) );
  XNOR2XL U332 ( .A(n205), .B(n206), .Y(n204) );
  XNOR2XL U333 ( .A(n207), .B(n208), .Y(n206) );
  XNOR2XL U334 ( .A(rxtx_buf[6]), .B(rxtx_buf[5]), .Y(n208) );
  XNOR2XL U335 ( .A(rxtx_buf[4]), .B(rxtx_buf[3]), .Y(n207) );
  XNOR2XL U336 ( .A(n209), .B(n210), .Y(n205) );
  XNOR2XL U337 ( .A(rxtx_buf[2]), .B(rxtx_buf[1]), .Y(n210) );
  XNOR2XL U338 ( .A(rxtx_buf[0]), .B(ff_idn), .Y(n209) );
  NAND2X1 U339 ( .A(n211), .B(n79), .Y(n160) );
  MUX2IX1 U340 ( .D0(n212), .D1(n213), .S(new_rx_sync_cnt[1]), .Y(N349) );
  AOI21X1 U341 ( .B(n214), .C(n161), .A(n215), .Y(n213) );
  NAND2X1 U342 ( .A(new_rx_sync_cnt[0]), .B(n214), .Y(n212) );
  MUX2X1 U343 ( .D0(n215), .D1(n214), .S(n161), .Y(N348) );
  INVX1 U344 ( .A(new_rx_sync_cnt[0]), .Y(n161) );
  AOI211X1 U345 ( .C(n216), .D(n217), .A(n117), .B(n214), .Y(n215) );
  OAI222XL U346 ( .A(n162), .B(n218), .C(n219), .D(n220), .E(n114), .F(n221), 
        .Y(n214) );
  INVX1 U347 ( .A(n195), .Y(n221) );
  OAI211X1 U348 ( .C(n180), .D(n526), .A(n198), .B(N331), .Y(n220) );
  NOR21XL U349 ( .B(n222), .A(n114), .Y(n526) );
  INVX1 U350 ( .A(n162), .Y(n180) );
  OAI2B11X1 U351 ( .D(n223), .C(n224), .A(n188), .B(n225), .Y(n219) );
  AOI32X1 U352 ( .A(n226), .B(n223), .C(n227), .D(ui_intv_cnt[6]), .E(n228), 
        .Y(n225) );
  INVX1 U353 ( .A(N338), .Y(n228) );
  AOI22AXL U354 ( .A(N336), .B(n187), .D(n229), .C(n230), .Y(n227) );
  NAND2X1 U355 ( .A(n14), .B(n231), .Y(n230) );
  OAI31XL U356 ( .A(n232), .B(n10), .C(n233), .D(n234), .Y(n229) );
  INVX1 U357 ( .A(n235), .Y(n234) );
  AOI211X1 U358 ( .C(n10), .D(n233), .A(n236), .B(n232), .Y(n235) );
  AOI22AXL U359 ( .A(n237), .B(ui_intv_cnt[0]), .D(N325), .C(ui_intv_cnt[1]), 
        .Y(n236) );
  AOI21X1 U360 ( .B(N325), .C(n86), .A(N324), .Y(n237) );
  NOR2X1 U361 ( .A(n231), .B(N141), .Y(n232) );
  INVX1 U362 ( .A(n361), .Y(n231) );
  AOI32X1 U363 ( .A(n226), .B(N328), .C(N142), .D(n7), .E(n238), .Y(n224) );
  INVX1 U364 ( .A(N337), .Y(n238) );
  NAND2X1 U365 ( .A(N337), .B(n88), .Y(n226) );
  NAND2X1 U366 ( .A(N338), .B(n87), .Y(n223) );
  NAND2X1 U367 ( .A(ff_chg), .B(n80), .Y(n162) );
  OAI21X1 U368 ( .B(n239), .C(n137), .A(n134), .Y(N261) );
  OAI211X1 U369 ( .C(n15), .D(n240), .A(n137), .B(n241), .Y(n134) );
  AOI21X1 U370 ( .B(n242), .C(n155), .A(n5), .Y(n241) );
  OAI22X1 U371 ( .A(n243), .B(n137), .C(n244), .D(n121), .Y(N260) );
  AOI22AXL U372 ( .A(n15), .B(n242), .D(n240), .C(n151), .Y(n244) );
  XNOR2XL U373 ( .A(n39), .B(ff_idn), .Y(n240) );
  XNOR2XL U374 ( .A(r_dat[7]), .B(n175), .Y(n242) );
  INVX1 U375 ( .A(n122), .Y(n137) );
  OAI211X1 U376 ( .C(n245), .D(n246), .A(n122), .B(n247), .Y(N22) );
  INVX1 U377 ( .A(n155), .Y(n151) );
  AOI31X1 U378 ( .A(n248), .B(n249), .C(n250), .D(n251), .Y(n164) );
  OAI31XL U379 ( .A(n252), .B(n253), .C(n254), .D(n255), .Y(n251) );
  NAND41X1 U380 ( .D(n256), .A(n257), .B(n258), .C(n259), .Y(n255) );
  AOI211X1 U381 ( .C(n260), .D(n18), .A(n261), .B(n262), .Y(n258) );
  INVX1 U382 ( .A(n263), .Y(n248) );
  NAND4X1 U383 ( .A(n264), .B(n265), .C(n266), .D(n267), .Y(N219) );
  NOR4XL U384 ( .A(n268), .B(n269), .C(n270), .D(n271), .Y(n267) );
  XNOR2XL U385 ( .A(ui_intv_cnt[0]), .B(n272), .Y(n271) );
  NAND21X1 U386 ( .B(n273), .A(r_tui[0]), .Y(n272) );
  AOI21X1 U387 ( .B(n92), .C(n80), .A(n274), .Y(n273) );
  XNOR2XL U388 ( .A(n275), .B(n87), .Y(n270) );
  ENOX1 U389 ( .A(n276), .B(n277), .C(adp_tx_ui_6_), .D(n274), .Y(n275) );
  XNOR2XL U390 ( .A(ui_intv_cnt[7]), .B(n278), .Y(n269) );
  AOI221XL U391 ( .A(n80), .B(rx_ui_1_2[6]), .C(n274), .D(adp_tx_ui_7_), .E(
        n117), .Y(n278) );
  XNOR2XL U392 ( .A(N142), .B(n279), .Y(n268) );
  AOI22X1 U393 ( .A(n274), .B(r_tui[4]), .C(n10), .D(n80), .Y(n279) );
  NOR2X1 U394 ( .A(n280), .B(n281), .Y(n266) );
  XNOR2XL U395 ( .A(n282), .B(n233), .Y(n281) );
  ENOX1 U396 ( .A(n276), .B(n172), .C(r_tui[2]), .D(n274), .Y(n282) );
  XNOR2XL U397 ( .A(N141), .B(n283), .Y(n280) );
  AOI22X1 U398 ( .A(n274), .B(r_tui[3]), .C(N325), .D(n80), .Y(n283) );
  XNOR2XL U399 ( .A(ui_intv_cnt[1]), .B(n284), .Y(n265) );
  ENOX1 U400 ( .A(n276), .B(n285), .C(r_tui[1]), .D(n274), .Y(n284) );
  XNOR2XL U401 ( .A(n286), .B(n88), .Y(n264) );
  AOI221XL U402 ( .A(n80), .B(rx_ui_1_2[4]), .C(n274), .D(adp_tx_ui_5_), .E(
        n117), .Y(n286) );
  NOR2X1 U403 ( .A(n2), .B(n117), .Y(n274) );
  NAND3X1 U404 ( .A(n168), .B(n167), .C(n169), .Y(N205) );
  INVX1 U405 ( .A(n171), .Y(n169) );
  OAI211X1 U406 ( .C(r_ctl[6]), .D(n114), .A(n155), .B(n247), .Y(n171) );
  OA21X1 U407 ( .B(n165), .C(n287), .A(n288), .Y(n247) );
  GEN2XL U408 ( .D(n260), .E(n289), .C(N363), .B(n290), .A(n291), .Y(n287) );
  AOI222XL U409 ( .A(n257), .B(n256), .C(n253), .D(n292), .E(n250), .F(n263), 
        .Y(n291) );
  OAI31XL U410 ( .A(n293), .B(n294), .C(n295), .D(n246), .Y(n263) );
  AOI21X1 U411 ( .B(N362), .C(n289), .A(N363), .Y(n295) );
  AOI21X1 U412 ( .B(N362), .C(n296), .A(n297), .Y(n294) );
  NAND2X1 U413 ( .A(n298), .B(n299), .Y(n250) );
  AOI21BBXL U414 ( .B(n300), .C(n301), .A(n302), .Y(n253) );
  AOI21X1 U415 ( .B(n303), .C(symb_cnt[2]), .A(symb_cnt[3]), .Y(n301) );
  AOI211X1 U416 ( .C(n304), .D(n305), .A(n306), .B(n307), .Y(n300) );
  OAI22X1 U417 ( .A(n303), .B(n308), .C(n303), .D(n297), .Y(n306) );
  NAND2X1 U418 ( .A(n243), .B(n296), .Y(n305) );
  OAI2B11X1 U419 ( .D(N419), .C(n293), .A(n309), .B(n246), .Y(n256) );
  NAND42X1 U420 ( .C(n310), .D(n311), .A(n312), .B(n313), .Y(n309) );
  NOR2X1 U421 ( .A(n262), .B(n261), .Y(n313) );
  NOR2X1 U422 ( .A(n297), .B(N418), .Y(n261) );
  NOR2X1 U423 ( .A(n308), .B(N419), .Y(n262) );
  OAI21X1 U424 ( .B(n18), .C(n260), .A(N160), .Y(n312) );
  INVX1 U425 ( .A(n243), .Y(n260) );
  AOI21X1 U426 ( .B(n296), .C(n243), .A(N418), .Y(n310) );
  OAI31XL U427 ( .A(n314), .B(n18), .C(n243), .D(n217), .Y(n290) );
  INVX1 U428 ( .A(N362), .Y(n243) );
  INVX1 U429 ( .A(n146), .Y(r_ctl[6]) );
  NAND32X1 U430 ( .B(n115), .C(n276), .A(ff_idn), .Y(n168) );
  AOI21X1 U431 ( .B(symb_cnt[3]), .C(n4), .A(n177), .Y(n115) );
  OAI211X1 U432 ( .C(n292), .D(n315), .A(n246), .B(n202), .Y(N1043) );
  ENOX1 U433 ( .A(n316), .B(n158), .C(n26), .D(n317), .Y(N1016) );
  INVX1 U434 ( .A(symb_cnt[6]), .Y(n158) );
  ENOX1 U435 ( .A(n316), .B(n318), .C(n27), .D(n317), .Y(N1015) );
  ENOX1 U436 ( .A(n316), .B(n319), .C(n28), .D(n317), .Y(N1014) );
  AO22X1 U437 ( .A(n11), .B(n320), .C(n29), .D(n317), .Y(N1013) );
  ENOX1 U438 ( .A(n316), .B(n308), .C(n30), .D(n317), .Y(N1012) );
  ENOX1 U439 ( .A(n316), .B(n297), .C(n31), .D(n317), .Y(N1011) );
  ENOX1 U440 ( .A(n316), .B(n296), .C(n32), .D(n317), .Y(N1010) );
  OAI221X1 U441 ( .A(n321), .B(n245), .C(n322), .D(n165), .E(n323), .Y(n317)
         );
  AOI31X1 U442 ( .A(ff_idn), .B(n324), .C(n325), .D(n326), .Y(n323) );
  OAI31XL U443 ( .A(n327), .B(n328), .C(n329), .D(n288), .Y(n326) );
  NAND32X1 U444 ( .B(n201), .C(n330), .A(n197), .Y(n288) );
  INVX1 U445 ( .A(n331), .Y(n325) );
  AOI222XL U446 ( .A(n332), .B(n333), .C(n330), .D(n334), .E(n292), .F(n335), 
        .Y(n322) );
  ENOX1 U447 ( .A(n254), .B(n299), .C(n249), .D(n257), .Y(n334) );
  INVX1 U448 ( .A(n211), .Y(n245) );
  NOR2X1 U449 ( .A(n336), .B(n276), .Y(n211) );
  INVX1 U450 ( .A(n337), .Y(n321) );
  AOI31X1 U451 ( .A(n332), .B(n333), .C(n165), .D(n320), .Y(n316) );
  OAI211X1 U452 ( .C(n196), .D(n338), .A(n339), .B(n340), .Y(n320) );
  AOI21X1 U453 ( .B(ff_idn), .C(n341), .A(n342), .Y(n340) );
  OAI21X1 U454 ( .B(n157), .C(n343), .A(n344), .Y(n341) );
  AOI32X1 U455 ( .A(n345), .B(n327), .C(n222), .D(n324), .E(n331), .Y(n344) );
  NAND4X1 U456 ( .A(n189), .B(n81), .C(n17), .D(ui_intv_cnt[6]), .Y(n331) );
  NOR43XL U457 ( .B(n86), .C(n233), .D(n346), .A(ui_intv_cnt[0]), .Y(n189) );
  NOR3XL U458 ( .A(N141), .B(n3), .C(ui_intv_cnt[5]), .Y(n346) );
  ENOX1 U459 ( .A(n176), .B(n173), .C(n343), .D(n347), .Y(n324) );
  NAND4X1 U460 ( .A(n17), .B(ui_intv_cnt[2]), .C(n348), .D(n349), .Y(n327) );
  NOR4XL U461 ( .A(ui_intv_cnt[7]), .B(ui_intv_cnt[6]), .C(ui_intv_cnt[1]), 
        .D(ui_intv_cnt[0]), .Y(n349) );
  NOR2X1 U462 ( .A(n167), .B(n350), .Y(n348) );
  XNOR2XL U463 ( .A(ui_intv_cnt[5]), .B(n66), .Y(n350) );
  INVX1 U464 ( .A(n328), .Y(n345) );
  NAND3X1 U465 ( .A(symb_cnt[6]), .B(n351), .C(symb_cnt[5]), .Y(n343) );
  NAND3X1 U466 ( .A(n333), .B(n319), .C(n308), .Y(n351) );
  INVX1 U467 ( .A(n347), .Y(n157) );
  AOI33X1 U468 ( .A(n352), .B(n197), .C(n201), .D(n337), .E(n336), .F(n80), 
        .Y(n339) );
  NAND4X1 U469 ( .A(n353), .B(n354), .C(n355), .D(n356), .Y(n336) );
  NOR4XL U470 ( .A(n167), .B(n357), .C(n358), .D(n359), .Y(n356) );
  XNOR2XL U471 ( .A(ui_intv_cnt[6]), .B(n360), .Y(n359) );
  XNOR2XL U472 ( .A(N142), .B(n361), .Y(n358) );
  XNOR2XL U473 ( .A(add_264_A_0_), .B(n78), .Y(n357) );
  INVX1 U474 ( .A(n285), .Y(add_264_A_0_) );
  NAND2X1 U475 ( .A(r_tui[1]), .B(n92), .Y(n285) );
  NOR3XL U476 ( .A(n362), .B(ui_intv_cnt[7]), .C(n363), .Y(n355) );
  XNOR2XL U477 ( .A(ui_intv_cnt[1]), .B(n172), .Y(n363) );
  MUX2IX1 U478 ( .D0(r_tui[2]), .D1(catch_sync[0]), .S(r_tui[7]), .Y(n172) );
  XNOR2XL U479 ( .A(gt_647_B_3_), .B(n88), .Y(n362) );
  XNOR2XL U480 ( .A(ui_intv_cnt[2]), .B(n16), .Y(n354) );
  XNOR2XL U481 ( .A(n14), .B(n10), .Y(n353) );
  OAI32X1 U482 ( .A(n218), .B(new_rx_sync_cnt[1]), .C(new_rx_sync_cnt[0]), .D(
        n365), .E(n366), .Y(n337) );
  NOR43XL U483 ( .B(rx_trans_8_chg), .C(n367), .D(ff_chg), .A(n368), .Y(n366)
         );
  OAI31XL U484 ( .A(n369), .B(ui_intv_cnt[6]), .C(n7), .D(n246), .Y(n368) );
  OAI21X1 U485 ( .B(rx_ui_1_2[6]), .C(n187), .A(n370), .Y(n369) );
  OAI22X1 U486 ( .A(N142), .B(n360), .C(n371), .D(n372), .Y(n370) );
  AOI211X1 U487 ( .C(n10), .D(n373), .A(n374), .B(n375), .Y(n372) );
  AOI21BBXL U488 ( .B(n373), .C(n10), .A(ui_intv_cnt[1]), .Y(n375) );
  OAI22X1 U489 ( .A(ui_intv_cnt[2]), .B(n361), .C(N141), .D(n277), .Y(n374) );
  NAND2X1 U490 ( .A(ui_intv_cnt[0]), .B(n364), .Y(n373) );
  MUX2IX1 U491 ( .D0(r_tui[3]), .D1(catch_sync[1]), .S(r_tui[7]), .Y(n364) );
  INVX1 U492 ( .A(r_tui[7]), .Y(n92) );
  MAJ3X1 U493 ( .A(n277), .B(n376), .C(N141), .Y(n371) );
  NOR2X1 U494 ( .A(rx_ui_1_2[4]), .B(n233), .Y(n376) );
  MUX2IX1 U495 ( .D0(adp_tx_ui_5_), .D1(catch_sync[3]), .S(r_tui[7]), .Y(n361)
         );
  MUX2IX1 U496 ( .D0(adp_tx_ui_6_), .D1(catch_sync[4]), .S(r_tui[7]), .Y(n277)
         );
  MUX2IX1 U497 ( .D0(adp_tx_ui_7_), .D1(catch_sync[5]), .S(r_tui[7]), .Y(n360)
         );
  OAI21X1 U498 ( .B(n377), .C(n378), .A(n379), .Y(n367) );
  OAI211X1 U499 ( .C(rx_ui_3_8[5]), .D(n88), .A(n380), .B(n381), .Y(n379) );
  AOI22AXL U500 ( .A(n382), .B(n383), .D(rx_ui_3_8[4]), .C(N142), .Y(n381) );
  NAND3X1 U501 ( .A(n384), .B(n385), .C(n386), .Y(n383) );
  AOI22AXL U502 ( .A(n387), .B(n388), .D(rx_ui_3_8[2]), .C(ui_intv_cnt[2]), 
        .Y(n386) );
  OAI21X1 U503 ( .B(n387), .C(n388), .A(ui_intv_cnt[1]), .Y(n384) );
  INVX1 U504 ( .A(rx_ui_3_8[1]), .Y(n388) );
  NAND2X1 U505 ( .A(rx_ui_3_8[0]), .B(n78), .Y(n387) );
  AOI32X1 U506 ( .A(n385), .B(n233), .C(rx_ui_3_8[2]), .D(rx_ui_3_8[3]), .E(
        n66), .Y(n382) );
  INVX1 U507 ( .A(ui_intv_cnt[2]), .Y(n233) );
  OR2X1 U508 ( .A(rx_ui_3_8[3]), .B(n66), .Y(n385) );
  INVX1 U509 ( .A(n378), .Y(n380) );
  OAI21X1 U510 ( .B(rx_ui_3_8[6]), .C(n87), .A(n188), .Y(n378) );
  AOI221XL U511 ( .A(rx_ui_3_8[5]), .B(n88), .C(rx_ui_3_8[6]), .D(n87), .E(
        n389), .Y(n377) );
  INVX1 U512 ( .A(n390), .Y(n389) );
  OAI211X1 U513 ( .C(n88), .D(rx_ui_3_8[5]), .A(rx_ui_3_8[4]), .B(n187), .Y(
        n390) );
  NAND4X1 U514 ( .A(n391), .B(n392), .C(n393), .D(n394), .Y(n201) );
  NOR4XL U515 ( .A(n395), .B(n396), .C(n397), .D(n398), .Y(n394) );
  XNOR2XL U516 ( .A(adp_tx_1_4[6]), .B(n87), .Y(n398) );
  XNOR2XL U517 ( .A(adp_tx_1_4[5]), .B(n88), .Y(n397) );
  XNOR2XL U518 ( .A(adp_tx_1_4[4]), .B(n187), .Y(n396) );
  XNOR2XL U519 ( .A(adp_tx_1_4[3]), .B(n66), .Y(n395) );
  NOR3XL U520 ( .A(n399), .B(ui_intv_cnt[7]), .C(n167), .Y(n393) );
  XNOR2XL U521 ( .A(adp_tx_1_4[0]), .B(n78), .Y(n399) );
  XNOR2XL U522 ( .A(ui_intv_cnt[1]), .B(adp_tx_1_4[1]), .Y(n392) );
  XNOR2XL U523 ( .A(ui_intv_cnt[2]), .B(adp_tx_1_4[2]), .Y(n391) );
  AOI21AX1 U524 ( .B(n330), .C(n197), .A(n400), .Y(n338) );
  AOI31X1 U525 ( .A(n332), .B(n308), .C(n289), .D(n292), .Y(n400) );
  INVX1 U526 ( .A(n352), .Y(n330) );
  OAI21X1 U527 ( .B(n239), .C(n217), .A(n401), .Y(n352) );
  OAI21X1 U528 ( .B(n260), .C(n296), .A(n402), .Y(n401) );
  OAI21X1 U529 ( .B(n239), .C(n314), .A(n217), .Y(n402) );
  INVX1 U530 ( .A(N159), .Y(n296) );
  INVX1 U531 ( .A(N363), .Y(n239) );
  NAND3X1 U532 ( .A(n403), .B(n404), .C(n405), .Y(N1009) );
  OA222X1 U533 ( .A(n406), .B(n407), .C(n408), .D(r_ctl[7]), .E(n252), .F(n409), .Y(n405) );
  OAI211X1 U534 ( .C(n407), .D(n406), .A(n410), .B(n411), .Y(N1008) );
  AOI32X1 U535 ( .A(r_ctl[0]), .B(n412), .C(r_ctl[1]), .D(n347), .E(r_ctl[5]), 
        .Y(n411) );
  NOR4XL U536 ( .A(n413), .B(fcp_state[0]), .C(fcp_state[1]), .D(fcp_state[3]), 
        .Y(n347) );
  OAI31XL U537 ( .A(n165), .B(r_ctl[7]), .C(n408), .D(n403), .Y(n412) );
  INVX1 U538 ( .A(n414), .Y(n403) );
  NOR2X1 U539 ( .A(n415), .B(n416), .Y(n408) );
  INVX1 U540 ( .A(n342), .Y(n410) );
  OAI32X1 U541 ( .A(n417), .B(n176), .C(n175), .D(n418), .E(n419), .Y(n342) );
  AOI21X1 U542 ( .B(fcp_state[2]), .C(n420), .A(n117), .Y(n176) );
  NOR4XL U543 ( .A(n421), .B(fcp_state[0]), .C(fcp_state[2]), .D(fcp_state[3]), 
        .Y(n117) );
  NAND31X1 U544 ( .C(n422), .A(n404), .B(n423), .Y(N1007) );
  AOI22AXL U545 ( .A(n424), .B(n425), .D(n329), .C(n328), .Y(n423) );
  OAI21X1 U546 ( .B(r_ctl[0]), .C(n426), .A(n140), .Y(n425) );
  NAND2X1 U547 ( .A(r_ctl[0]), .B(n426), .Y(n140) );
  GEN2XL U548 ( .D(n409), .E(n292), .C(n415), .B(n163), .A(n414), .Y(n424) );
  OA222X1 U549 ( .A(n427), .B(n298), .C(n418), .D(n419), .E(n428), .F(n299), 
        .Y(n404) );
  NAND3X1 U550 ( .A(n365), .B(n80), .C(ff_idn), .Y(n419) );
  INVX1 U551 ( .A(n216), .Y(n365) );
  NOR3XL U552 ( .A(n165), .B(n429), .C(n315), .Y(n427) );
  OAI211X1 U553 ( .C(n328), .D(n329), .A(n430), .B(n431), .Y(N1006) );
  AOI221XL U554 ( .A(n292), .B(n432), .C(n433), .D(n434), .E(n422), .Y(n431)
         );
  NAND2X1 U555 ( .A(n435), .B(n436), .Y(n422) );
  NAND4X1 U556 ( .A(n222), .B(n198), .C(n18), .D(n175), .Y(n436) );
  OAI21X1 U557 ( .B(n418), .C(n216), .A(n80), .Y(n435) );
  INVX1 U558 ( .A(n218), .Y(n418) );
  NAND4X1 U559 ( .A(n18), .B(n437), .C(symb_cnt[3]), .D(n297), .Y(n218) );
  INVX1 U560 ( .A(n409), .Y(n432) );
  NOR3XL U561 ( .A(n246), .B(n165), .C(n335), .Y(n409) );
  INVX1 U562 ( .A(n252), .Y(n292) );
  AOI32X1 U563 ( .A(r_ctl[4]), .B(n195), .C(n438), .D(n439), .E(n426), .Y(n430) );
  INVX1 U564 ( .A(r_ctl[1]), .Y(n426) );
  GEN2XL U565 ( .D(n415), .E(n196), .C(n416), .B(n163), .A(n414), .Y(n439) );
  OAI32X1 U566 ( .A(n440), .B(n438), .C(n155), .D(r_ctl[7]), .E(n441), .Y(n414) );
  AOI22X1 U567 ( .A(n428), .B(n433), .C(n407), .D(n257), .Y(n441) );
  NOR2X1 U568 ( .A(n249), .B(n165), .Y(n407) );
  GEN2XL U569 ( .D(n260), .E(n297), .C(n442), .B(n437), .A(n216), .Y(n249) );
  NAND2X1 U570 ( .A(n246), .B(n315), .Y(n216) );
  OA21X1 U571 ( .B(n443), .C(N362), .A(N363), .Y(n442) );
  INVX1 U572 ( .A(n299), .Y(n433) );
  INVX1 U573 ( .A(n434), .Y(n428) );
  NAND2X1 U574 ( .A(n196), .B(n254), .Y(n434) );
  GEN3XL U575 ( .F(N362), .G(N159), .E(N160), .D(n444), .C(symb_cnt[2]), .B(
        symb_cnt[3]), .A(n302), .Y(n254) );
  OAI21BBX1 U576 ( .A(symb_cnt[3]), .B(n303), .C(n259), .Y(n302) );
  NOR2X1 U577 ( .A(n304), .B(N362), .Y(n303) );
  INVX1 U578 ( .A(n445), .Y(n304) );
  NAND2X1 U579 ( .A(n445), .B(n443), .Y(n444) );
  XNOR2XL U580 ( .A(N363), .B(N362), .Y(n445) );
  NAND2X1 U581 ( .A(n195), .B(r_wr[3]), .Y(n155) );
  INVX1 U582 ( .A(r_ctl[4]), .Y(n440) );
  INVX1 U583 ( .A(r_ctl[7]), .Y(n163) );
  NOR3XL U584 ( .A(n246), .B(n252), .C(n335), .Y(n416) );
  NAND2X1 U585 ( .A(n307), .B(symb_cnt[2]), .Y(n335) );
  INVX1 U586 ( .A(n443), .Y(n307) );
  NAND2X1 U587 ( .A(N159), .B(N160), .Y(n443) );
  INVX1 U588 ( .A(n165), .Y(n196) );
  NOR4XL U589 ( .A(n450), .B(n451), .C(n452), .D(n453), .Y(n449) );
  XNOR2XL U590 ( .A(n188), .B(adp_tx_ui_7_), .Y(n453) );
  INVX1 U591 ( .A(ui_intv_cnt[7]), .Y(n188) );
  XNOR2XL U592 ( .A(n87), .B(adp_tx_ui_6_), .Y(n452) );
  INVX1 U593 ( .A(ui_intv_cnt[6]), .Y(n87) );
  XNOR2XL U594 ( .A(n88), .B(adp_tx_ui_5_), .Y(n451) );
  XNOR2XL U595 ( .A(n187), .B(r_tui[4]), .Y(n450) );
  INVX1 U596 ( .A(N142), .Y(n187) );
  NOR3XL U597 ( .A(n454), .B(n167), .C(n455), .Y(n448) );
  XNOR2XL U598 ( .A(r_tui[1]), .B(n86), .Y(n455) );
  INVX1 U599 ( .A(ui_intv_cnt[1]), .Y(n86) );
  INVX1 U600 ( .A(n81), .Y(n167) );
  NOR42XL U601 ( .C(us_cnt[3]), .D(n192), .A(n195), .B(us_cnt[2]), .Y(n81) );
  INVX1 U602 ( .A(n194), .Y(n192) );
  NAND2X1 U603 ( .A(us_cnt[1]), .B(us_cnt[0]), .Y(n194) );
  XNOR2XL U604 ( .A(n78), .B(r_tui[0]), .Y(n454) );
  INVX1 U605 ( .A(ui_intv_cnt[0]), .Y(n78) );
  XNOR2XL U606 ( .A(ui_intv_cnt[2]), .B(r_tui[2]), .Y(n447) );
  XNOR2XL U607 ( .A(N141), .B(r_tui[3]), .Y(n446) );
  AND2X1 U608 ( .A(n79), .B(n332), .Y(n415) );
  INVX1 U609 ( .A(n298), .Y(n332) );
  NOR2X1 U610 ( .A(n315), .B(n333), .Y(n79) );
  NAND2X1 U611 ( .A(n437), .B(n289), .Y(n315) );
  INVX1 U612 ( .A(n293), .Y(n437) );
  NAND2X1 U613 ( .A(n259), .B(n308), .Y(n293) );
  NOR3XL U614 ( .A(n114), .B(n18), .C(n217), .Y(n438) );
  INVX1 U615 ( .A(n198), .Y(n217) );
  NOR2X1 U616 ( .A(n314), .B(N160), .Y(n198) );
  INVX1 U617 ( .A(ff_chg), .Y(n114) );
  NOR4XL U618 ( .A(fcp_state[0]), .B(fcp_state[1]), .C(fcp_state[2]), .D(
        fcp_state[3]), .Y(n195) );
  NAND2X1 U619 ( .A(n222), .B(ff_idn), .Y(n329) );
  NOR32XL U620 ( .B(n421), .C(n456), .A(fcp_state[3]), .Y(n222) );
  NOR3XL U621 ( .A(n297), .B(n18), .C(n314), .Y(n328) );
  NAND2X1 U622 ( .A(n429), .B(n308), .Y(n314) );
  INVX1 U623 ( .A(n246), .Y(n429) );
  INVX1 U624 ( .A(N160), .Y(n297) );
  NAND4X1 U625 ( .A(n276), .B(n146), .C(n457), .D(n458), .Y(N1005) );
  AOI211X1 U626 ( .C(ff_chg), .D(n177), .A(n175), .B(n421), .Y(n458) );
  INVX1 U627 ( .A(ff_idn), .Y(n175) );
  OAI21X1 U628 ( .B(n333), .C(n308), .A(n259), .Y(n177) );
  AOI21X1 U629 ( .B(fcp_state[2]), .C(n459), .A(n173), .Y(n457) );
  INVX1 U630 ( .A(n417), .Y(n173) );
  OAI31XL U631 ( .A(n460), .B(symb_cnt[6]), .C(symb_cnt[5]), .D(n311), .Y(n417) );
  INVX1 U632 ( .A(n259), .Y(n311) );
  NOR2X1 U633 ( .A(n159), .B(symb_cnt[6]), .Y(n259) );
  NAND2X1 U634 ( .A(n318), .B(n319), .Y(n159) );
  INVX1 U635 ( .A(symb_cnt[4]), .Y(n319) );
  INVX1 U636 ( .A(symb_cnt[5]), .Y(n318) );
  OAI21X1 U637 ( .B(n289), .C(n308), .A(n333), .Y(n460) );
  INVX1 U638 ( .A(symb_cnt[3]), .Y(n333) );
  NOR2X1 U639 ( .A(N160), .B(N159), .Y(n289) );
  NOR2X1 U640 ( .A(n197), .B(n202), .Y(n146) );
  NAND2X1 U641 ( .A(n298), .B(n252), .Y(n202) );
  NAND3X1 U642 ( .A(n456), .B(n421), .C(fcp_state[3]), .Y(n252) );
  NAND2X1 U643 ( .A(n420), .B(n413), .Y(n298) );
  NOR2X1 U644 ( .A(n459), .B(n421), .Y(n420) );
  NAND2X1 U645 ( .A(n299), .B(n406), .Y(n197) );
  INVX1 U646 ( .A(n257), .Y(n406) );
  NOR3XL U647 ( .A(n459), .B(fcp_state[1]), .C(n413), .Y(n257) );
  NAND21X1 U648 ( .B(fcp_state[0]), .A(fcp_state[3]), .Y(n459) );
  NAND3X1 U649 ( .A(fcp_state[1]), .B(n456), .C(fcp_state[3]), .Y(n299) );
  NAND32X1 U650 ( .B(fcp_state[3]), .C(n421), .A(n456), .Y(n276) );
  AND2X1 U651 ( .A(fcp_state[0]), .B(n413), .Y(n456) );
  INVX1 U652 ( .A(fcp_state[2]), .Y(n413) );
  INVX1 U653 ( .A(fcp_state[1]), .Y(n421) );
endmodule


module fcpegn_a0_DW01_inc_2 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  XOR2X1 U1 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module fcpegn_a0_DW01_inc_1 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [6:2] carry;

  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(SUM[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
endmodule


module fcpegn_a0_DW01_inc_0 ( A, SUM );
  input [6:0] A;
  output [6:0] SUM;

  wire   [6:2] carry;

  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  XOR2X1 U1 ( .A(carry[6]), .B(A[6]), .Y(SUM[6]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_fcpegn_a0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_fcpegn_a0_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_fcpegn_a0_3 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_fcpegn_a0_4 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_fcpegn_a0_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_2 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net9515;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_2 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9515), .TE(1'b0) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net9515), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net9515), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net9515), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net9515), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net9515), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net9515), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net9515), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net9515), .XR(arstz), .Q(rdat[4]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_3 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net9533;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_3 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9533), .TE(1'b0) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net9533), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net9533), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net9533), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net9533), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net9533), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net9533), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net9533), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net9533), .XR(arstz), .Q(rdat[4]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_3 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_4 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net9551;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_4 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9551), .TE(1'b0) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net9551), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net9551), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net9551), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net9551), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net9551), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net9551), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net9551), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net9551), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_4 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glsta_a0_0 ( clk, arstz, rst0, set2, clr1, rdat, irq );
  input [7:0] set2;
  input [7:0] clr1;
  output [7:0] rdat;
  output [7:0] irq;
  input clk, arstz, rst0;
  wire   upd_r, n17, n18, n19, n20, n21, n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16;
  wire   [7:0] wd_r;

  glreg_WIDTH8_0 u0 ( .clk(clk), .arstz(arstz), .we(upd_r), .wdat(wd_r), 
        .rdat(rdat) );
  NOR4XL U2 ( .A(clr1[7]), .B(clr1[6]), .C(clr1[5]), .D(clr1[4]), .Y(n18) );
  INVX1 U3 ( .A(set2[4]), .Y(n2) );
  INVX1 U4 ( .A(set2[0]), .Y(n3) );
  INVX1 U5 ( .A(set2[1]), .Y(n1) );
  INVX1 U6 ( .A(set2[2]), .Y(n7) );
  NAND3X1 U7 ( .A(n6), .B(n4), .C(n16), .Y(n21) );
  INVX1 U8 ( .A(set2[6]), .Y(n6) );
  INVX1 U9 ( .A(set2[3]), .Y(n5) );
  NAND4X1 U10 ( .A(n17), .B(n18), .C(n19), .D(n20), .Y(upd_r) );
  NOR4XL U11 ( .A(set2[2]), .B(set2[1]), .C(set2[0]), .D(rst0), .Y(n19) );
  NOR3XL U12 ( .A(n21), .B(set2[4]), .C(set2[3]), .Y(n20) );
  NOR4XL U13 ( .A(clr1[3]), .B(clr1[2]), .C(clr1[1]), .D(clr1[0]), .Y(n17) );
  AOI211X1 U14 ( .C(n3), .D(n15), .A(rst0), .B(clr1[0]), .Y(wd_r[0]) );
  INVX1 U15 ( .A(rdat[0]), .Y(n15) );
  AOI211X1 U16 ( .C(n1), .D(n14), .A(rst0), .B(clr1[1]), .Y(wd_r[1]) );
  INVX1 U17 ( .A(rdat[1]), .Y(n14) );
  AOI211X1 U18 ( .C(n7), .D(n13), .A(rst0), .B(clr1[2]), .Y(wd_r[2]) );
  INVX1 U19 ( .A(rdat[2]), .Y(n13) );
  AOI211X1 U20 ( .C(n5), .D(n12), .A(rst0), .B(clr1[3]), .Y(wd_r[3]) );
  INVX1 U21 ( .A(rdat[3]), .Y(n12) );
  AOI211X1 U22 ( .C(n2), .D(n11), .A(rst0), .B(clr1[4]), .Y(wd_r[4]) );
  INVX1 U23 ( .A(rdat[4]), .Y(n11) );
  AOI211X1 U24 ( .C(n16), .D(n10), .A(rst0), .B(clr1[5]), .Y(wd_r[5]) );
  INVX1 U25 ( .A(rdat[5]), .Y(n10) );
  AOI211X1 U26 ( .C(n6), .D(n9), .A(rst0), .B(clr1[6]), .Y(wd_r[6]) );
  INVX1 U27 ( .A(rdat[6]), .Y(n9) );
  AOI211X1 U28 ( .C(n4), .D(n8), .A(rst0), .B(clr1[7]), .Y(wd_r[7]) );
  INVX1 U29 ( .A(rdat[7]), .Y(n8) );
  NOR2X1 U30 ( .A(rdat[6]), .B(n6), .Y(irq[6]) );
  NOR2X1 U31 ( .A(rdat[7]), .B(n4), .Y(irq[7]) );
  INVX1 U32 ( .A(set2[7]), .Y(n4) );
  NOR2X1 U33 ( .A(rdat[5]), .B(n16), .Y(irq[5]) );
  NOR2X1 U34 ( .A(rdat[4]), .B(n2), .Y(irq[4]) );
  NOR2X1 U35 ( .A(rdat[1]), .B(n1), .Y(irq[1]) );
  NOR2X1 U36 ( .A(rdat[0]), .B(n3), .Y(irq[0]) );
  NOR2X1 U37 ( .A(rdat[2]), .B(n7), .Y(irq[2]) );
  NOR2X1 U38 ( .A(rdat[3]), .B(n5), .Y(irq[3]) );
  INVX1 U39 ( .A(set2[5]), .Y(n16) );
endmodule


module glreg_WIDTH8_0 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net9569;

  SNPS_CLOCK_GATE_HIGH_glreg_WIDTH8_0 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9569), .TE(1'b0) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net9569), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net9569), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net9569), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net9569), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net9569), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net9569), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net9569), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net9569), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_WIDTH8_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_8_00000000 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net9587;

  SNPS_CLOCK_GATE_HIGH_glreg_8_00000000 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9587), .TE(1'b0) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net9587), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net9587), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net9587), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net9587), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net9587), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net9587), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net9587), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net9587), .XR(arstz), .Q(rdat[6]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_8_00000000 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module dpdmacc_a0 ( dp_comp, dm_comp, id_comp, r_re_0, r_wr_1, r_wdat, r_acc, 
        r_dpdmsta, r_dm, r_dmchg, r_int, clk, rstz );
  input [7:0] r_wdat;
  output [7:0] r_acc;
  output [7:0] r_dpdmsta;
  input dp_comp, dm_comp, id_comp, r_re_0, r_wr_1, clk, rstz;
  output r_dm, r_dmchg, r_int;
  wire   dp_chg, dp_rise, dm_fall, dp_active_acc, dp_inacti_acc, dm_active_acc,
         dm_inacti_acc, upd00, N12, N15, N16, N17, N18, N19, N22, N23, N24,
         N25, n21, n22, n23, n24, n25, n26, N34, N35, n1, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20;
  wire   [7:0] wd00;

  ff_sync_2 u0_dpsync ( .i_org(dp_comp), .o_dbc(r_dpdmsta[6]), .o_chg(dp_chg), 
        .clk(clk), .rstz(n4) );
  ff_sync_1 u0_dmsync ( .i_org(dm_comp), .o_dbc(r_dpdmsta[7]), .o_chg(r_dmchg), 
        .clk(clk), .rstz(n4) );
  ff_sync_0 u0_idsync ( .i_org(id_comp), .o_dbc(r_dpdmsta[5]), .o_chg(), .clk(
        clk), .rstz(n5) );
  filter150us_a0_1 u0_dpfltr ( .active_hit(dp_active_acc), .inacti_hit(
        dp_inacti_acc), .start_edge(dp_rise), .any_edge(dp_chg), .clk(clk), 
        .rstz(n5) );
  filter150us_a0_0 u0_dmfltr ( .active_hit(dm_active_acc), .inacti_hit(
        dm_inacti_acc), .start_edge(dm_fall), .any_edge(r_dmchg), .clk(clk), 
        .rstz(n5) );
  glreg_a0_5 u0_accmltr ( .clk(clk), .arstz(n3), .we(upd00), .wdat(wd00), 
        .rdat(r_acc) );
  glreg_WIDTH5_0 u0_dpdmsta ( .clk(clk), .arstz(n4), .we(r_wr_1), .wdat(
        r_wdat[4:0]), .rdat(r_dpdmsta[4:0]) );
  INVX1 U3 ( .A(r_re_0), .Y(n1) );
  INVX1 U4 ( .A(n8), .Y(r_dm) );
  INVX1 U5 ( .A(n6), .Y(n4) );
  INVX1 U6 ( .A(n6), .Y(n3) );
  INVX1 U7 ( .A(n6), .Y(n5) );
  INVX1 U8 ( .A(rstz), .Y(n6) );
  NAND2X1 U9 ( .A(n23), .B(n1), .Y(upd00) );
  INVX1 U10 ( .A(r_re_0), .Y(n9) );
  NOR2X1 U11 ( .A(n7), .B(n11), .Y(n23) );
  NOR21XL U12 ( .B(r_dmchg), .A(n8), .Y(dm_fall) );
  INVX1 U13 ( .A(n22), .Y(n11) );
  INVX1 U14 ( .A(n21), .Y(n7) );
  OAI21X1 U15 ( .B(n23), .C(n9), .A(n24), .Y(r_int) );
  AOI33X1 U16 ( .A(n7), .B(n13), .C(n25), .D(n11), .E(n14), .F(n26), .Y(n24)
         );
  INVX1 U17 ( .A(r_acc[0]), .Y(n14) );
  AND2X1 U18 ( .A(N23), .B(n9), .Y(wd00[1]) );
  XNOR2XL U19 ( .A(r_acc[1]), .B(n20), .Y(N23) );
  AND2X1 U20 ( .A(N24), .B(n9), .Y(wd00[2]) );
  XOR2X1 U21 ( .A(n19), .B(r_acc[2]), .Y(N24) );
  NOR21XL U22 ( .B(r_acc[1]), .A(n20), .Y(n19) );
  AND2X1 U23 ( .A(N25), .B(n9), .Y(wd00[3]) );
  XNOR2XL U24 ( .A(r_acc[3]), .B(n18), .Y(N25) );
  NAND4X1 U25 ( .A(r_acc[2]), .B(r_acc[1]), .C(N34), .D(r_acc[0]), .Y(n18) );
  AND2X1 U26 ( .A(N16), .B(n9), .Y(wd00[5]) );
  XNOR2XL U27 ( .A(r_acc[5]), .B(n17), .Y(N16) );
  AND2X1 U28 ( .A(N17), .B(n9), .Y(wd00[6]) );
  XOR2X1 U29 ( .A(n16), .B(r_acc[6]), .Y(N17) );
  NOR21XL U30 ( .B(r_acc[5]), .A(n17), .Y(n16) );
  AND2X1 U31 ( .A(N18), .B(n9), .Y(wd00[7]) );
  XNOR2XL U32 ( .A(r_acc[7]), .B(n15), .Y(N18) );
  NAND4X1 U33 ( .A(r_acc[6]), .B(r_acc[5]), .C(N35), .D(r_acc[4]), .Y(n15) );
  ENOX1 U34 ( .A(n22), .B(n9), .C(N22), .D(n9), .Y(wd00[0]) );
  XOR2X1 U35 ( .A(N34), .B(r_acc[0]), .Y(N22) );
  ENOX1 U36 ( .A(n21), .B(n1), .C(N15), .D(n9), .Y(wd00[4]) );
  XOR2X1 U37 ( .A(N35), .B(r_acc[4]), .Y(N15) );
  AOI32X1 U38 ( .A(n10), .B(n8), .C(dm_active_acc), .D(r_dpdmsta[1]), .E(
        dm_inacti_acc), .Y(n21) );
  INVX1 U39 ( .A(r_dpdmsta[1]), .Y(n10) );
  AOI32X1 U40 ( .A(dp_active_acc), .B(n12), .C(r_dpdmsta[6]), .D(r_dpdmsta[0]), 
        .E(dp_inacti_acc), .Y(n22) );
  INVX1 U41 ( .A(r_dpdmsta[0]), .Y(n12) );
  NOR21XL U42 ( .B(dp_chg), .A(r_dpdmsta[6]), .Y(dp_rise) );
  INVX1 U43 ( .A(r_dpdmsta[7]), .Y(n8) );
  AND2X1 U44 ( .A(N19), .B(n11), .Y(N34) );
  NAND4X1 U45 ( .A(r_acc[3]), .B(r_acc[2]), .C(r_acc[1]), .D(r_acc[0]), .Y(N19) );
  AND2X1 U46 ( .A(N12), .B(n7), .Y(N35) );
  NAND4X1 U47 ( .A(r_acc[7]), .B(r_acc[6]), .C(r_acc[5]), .D(r_acc[4]), .Y(N12) );
  NAND2X1 U48 ( .A(N34), .B(r_acc[0]), .Y(n20) );
  NAND2X1 U49 ( .A(N35), .B(r_acc[4]), .Y(n17) );
  NOR3XL U50 ( .A(r_acc[1]), .B(r_acc[3]), .C(r_acc[2]), .Y(n26) );
  NOR3XL U51 ( .A(r_acc[5]), .B(r_acc[7]), .C(r_acc[6]), .Y(n25) );
  INVX1 U52 ( .A(r_acc[4]), .Y(n13) );
endmodule


module glreg_WIDTH5_0 ( clk, arstz, we, wdat, rdat );
  input [4:0] wdat;
  output [4:0] rdat;
  input clk, arstz, we;
  wire   net9605;

  SNPS_CLOCK_GATE_HIGH_glreg_WIDTH5_0 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9605), .TE(1'b0) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net9605), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net9605), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net9605), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net9605), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net9605), .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_WIDTH5_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_5 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net9623;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_5 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9623), .TE(1'b0) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net9623), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net9623), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net9623), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net9623), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net9623), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net9623), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net9623), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net9623), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_5 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module filter150us_a0_0 ( active_hit, inacti_hit, start_edge, any_edge, clk, 
        rstz );
  input start_edge, any_edge, clk, rstz;
  output active_hit, inacti_hit;
  wire   N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24, N25,
         N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, net9641, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16;
  wire   [11:0] dbcnt;

  SNPS_CLOCK_GATE_HIGH_filter150us_a0_0 clk_gate_dbcnt_reg ( .CLK(clk), .EN(
        N24), .ENCLK(net9641), .TE(1'b0) );
  filter150us_a0_0_DW01_inc_0 add_76 ( .A(dbcnt), .SUM({N23, N22, N21, N20, 
        N19, N18, N17, N16, N15, N14, N13, N12}) );
  DFFRQX1 dbcnt_reg_11_ ( .D(N36), .C(net9641), .XR(n2), .Q(dbcnt[11]) );
  DFFRQX1 dbcnt_reg_1_ ( .D(N26), .C(net9641), .XR(rstz), .Q(dbcnt[1]) );
  DFFRQX1 dbcnt_reg_9_ ( .D(N34), .C(net9641), .XR(n2), .Q(dbcnt[9]) );
  DFFRQX1 dbcnt_reg_2_ ( .D(N27), .C(net9641), .XR(rstz), .Q(dbcnt[2]) );
  DFFRQX1 dbcnt_reg_8_ ( .D(N33), .C(net9641), .XR(n2), .Q(dbcnt[8]) );
  DFFRQX1 dbcnt_reg_10_ ( .D(N35), .C(net9641), .XR(n2), .Q(dbcnt[10]) );
  DFFRQX1 dbcnt_reg_0_ ( .D(N25), .C(net9641), .XR(n2), .Q(dbcnt[0]) );
  DFFRQX1 dbcnt_reg_6_ ( .D(N31), .C(net9641), .XR(n2), .Q(dbcnt[6]) );
  DFFRQX1 dbcnt_reg_5_ ( .D(N30), .C(net9641), .XR(n2), .Q(dbcnt[5]) );
  DFFRQX1 dbcnt_reg_7_ ( .D(N32), .C(net9641), .XR(n2), .Q(dbcnt[7]) );
  DFFRQX1 dbcnt_reg_3_ ( .D(N28), .C(net9641), .XR(n2), .Q(dbcnt[3]) );
  DFFRQX1 dbcnt_reg_4_ ( .D(N29), .C(net9641), .XR(n2), .Q(dbcnt[4]) );
  BUFX3 U3 ( .A(n11), .Y(n1) );
  INVX1 U4 ( .A(n3), .Y(n2) );
  INVX1 U5 ( .A(rstz), .Y(n3) );
  NOR3XL U6 ( .A(n13), .B(any_edge), .C(n14), .Y(n11) );
  AOI211X1 U7 ( .C(n4), .D(n5), .A(n6), .B(start_edge), .Y(inacti_hit) );
  INVX1 U8 ( .A(any_edge), .Y(n6) );
  AO21X1 U9 ( .B(n7), .C(n8), .A(n9), .Y(n5) );
  NOR4XL U10 ( .A(dbcnt[11]), .B(n10), .C(n9), .D(n7), .Y(active_hit) );
  NAND3X1 U11 ( .A(dbcnt[1]), .B(dbcnt[0]), .C(dbcnt[2]), .Y(n7) );
  AND2X1 U12 ( .A(N23), .B(n1), .Y(N36) );
  AND2X1 U13 ( .A(N22), .B(n1), .Y(N35) );
  AND2X1 U14 ( .A(N21), .B(n1), .Y(N34) );
  AND2X1 U15 ( .A(N20), .B(n1), .Y(N33) );
  AND2X1 U16 ( .A(N19), .B(n11), .Y(N32) );
  AND2X1 U17 ( .A(N18), .B(n11), .Y(N31) );
  AND2X1 U18 ( .A(N17), .B(n11), .Y(N30) );
  AND2X1 U19 ( .A(N16), .B(n11), .Y(N29) );
  AND2X1 U20 ( .A(N15), .B(n11), .Y(N28) );
  AND2X1 U21 ( .A(N14), .B(n11), .Y(N27) );
  AND2X1 U22 ( .A(N13), .B(n11), .Y(N26) );
  OAI21BBX1 U23 ( .A(N12), .B(n11), .C(n12), .Y(N25) );
  OAI21X1 U24 ( .B(n13), .C(n14), .A(any_edge), .Y(n12) );
  OR2X1 U25 ( .A(n11), .B(any_edge), .Y(N24) );
  OAI21X1 U26 ( .B(n8), .C(n9), .A(n4), .Y(n14) );
  INVX1 U27 ( .A(dbcnt[11]), .Y(n4) );
  NAND3X1 U28 ( .A(dbcnt[8]), .B(dbcnt[10]), .C(dbcnt[9]), .Y(n9) );
  NOR42XL U29 ( .C(n8), .D(n15), .A(dbcnt[0]), .B(dbcnt[10]), .Y(n13) );
  NOR4XL U30 ( .A(dbcnt[9]), .B(dbcnt[8]), .C(dbcnt[2]), .D(dbcnt[1]), .Y(n15)
         );
  INVX1 U31 ( .A(n10), .Y(n8) );
  NAND32X1 U32 ( .B(dbcnt[4]), .C(dbcnt[3]), .A(n16), .Y(n10) );
  NOR3XL U33 ( .A(dbcnt[5]), .B(dbcnt[7]), .C(dbcnt[6]), .Y(n16) );
endmodule


module filter150us_a0_0_DW01_inc_0 ( A, SUM );
  input [11:0] A;
  output [11:0] SUM;

  wire   [11:2] carry;

  HAD1X1 U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .SO(SUM[10]) );
  HAD1X1 U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .SO(SUM[9]) );
  HAD1X1 U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .SO(SUM[8]) );
  HAD1X1 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .SO(SUM[7]) );
  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  XOR2X1 U1 ( .A(carry[11]), .B(A[11]), .Y(SUM[11]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_filter150us_a0_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module filter150us_a0_1 ( active_hit, inacti_hit, start_edge, any_edge, clk, 
        rstz );
  input start_edge, any_edge, clk, rstz;
  output active_hit, inacti_hit;
  wire   N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24, N25,
         N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, net9659, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16;
  wire   [11:0] dbcnt;

  SNPS_CLOCK_GATE_HIGH_filter150us_a0_1 clk_gate_dbcnt_reg ( .CLK(clk), .EN(
        N24), .ENCLK(net9659), .TE(1'b0) );
  filter150us_a0_1_DW01_inc_0 add_76 ( .A(dbcnt), .SUM({N23, N22, N21, N20, 
        N19, N18, N17, N16, N15, N14, N13, N12}) );
  DFFRQX1 dbcnt_reg_4_ ( .D(N29), .C(net9659), .XR(n2), .Q(dbcnt[4]) );
  DFFRQX1 dbcnt_reg_11_ ( .D(N36), .C(net9659), .XR(n2), .Q(dbcnt[11]) );
  DFFRQX1 dbcnt_reg_1_ ( .D(N26), .C(net9659), .XR(rstz), .Q(dbcnt[1]) );
  DFFRQX1 dbcnt_reg_9_ ( .D(N34), .C(net9659), .XR(n2), .Q(dbcnt[9]) );
  DFFRQX1 dbcnt_reg_2_ ( .D(N27), .C(net9659), .XR(rstz), .Q(dbcnt[2]) );
  DFFRQX1 dbcnt_reg_8_ ( .D(N33), .C(net9659), .XR(n2), .Q(dbcnt[8]) );
  DFFRQX1 dbcnt_reg_10_ ( .D(N35), .C(net9659), .XR(n2), .Q(dbcnt[10]) );
  DFFRQX1 dbcnt_reg_0_ ( .D(N25), .C(net9659), .XR(n2), .Q(dbcnt[0]) );
  DFFRQX1 dbcnt_reg_6_ ( .D(N31), .C(net9659), .XR(n2), .Q(dbcnt[6]) );
  DFFRQX1 dbcnt_reg_5_ ( .D(N30), .C(net9659), .XR(n2), .Q(dbcnt[5]) );
  DFFRQX1 dbcnt_reg_7_ ( .D(N32), .C(net9659), .XR(n2), .Q(dbcnt[7]) );
  DFFRQX1 dbcnt_reg_3_ ( .D(N28), .C(net9659), .XR(n2), .Q(dbcnt[3]) );
  BUFX3 U3 ( .A(n11), .Y(n1) );
  INVX1 U4 ( .A(n3), .Y(n2) );
  INVX1 U5 ( .A(rstz), .Y(n3) );
  NOR3XL U6 ( .A(n13), .B(any_edge), .C(n14), .Y(n11) );
  AOI211X1 U7 ( .C(n4), .D(n5), .A(n6), .B(start_edge), .Y(inacti_hit) );
  INVX1 U8 ( .A(any_edge), .Y(n6) );
  AO21X1 U9 ( .B(n7), .C(n8), .A(n9), .Y(n5) );
  NOR4XL U10 ( .A(dbcnt[11]), .B(n10), .C(n9), .D(n7), .Y(active_hit) );
  NAND3X1 U11 ( .A(dbcnt[1]), .B(dbcnt[0]), .C(dbcnt[2]), .Y(n7) );
  AND2X1 U12 ( .A(N23), .B(n1), .Y(N36) );
  AND2X1 U13 ( .A(N22), .B(n1), .Y(N35) );
  AND2X1 U14 ( .A(N21), .B(n1), .Y(N34) );
  AND2X1 U15 ( .A(N20), .B(n1), .Y(N33) );
  AND2X1 U16 ( .A(N19), .B(n11), .Y(N32) );
  AND2X1 U17 ( .A(N18), .B(n11), .Y(N31) );
  AND2X1 U18 ( .A(N17), .B(n11), .Y(N30) );
  AND2X1 U19 ( .A(N16), .B(n11), .Y(N29) );
  AND2X1 U20 ( .A(N15), .B(n11), .Y(N28) );
  AND2X1 U21 ( .A(N14), .B(n11), .Y(N27) );
  AND2X1 U22 ( .A(N13), .B(n11), .Y(N26) );
  OAI21BBX1 U23 ( .A(N12), .B(n11), .C(n12), .Y(N25) );
  OAI21X1 U24 ( .B(n13), .C(n14), .A(any_edge), .Y(n12) );
  OR2X1 U25 ( .A(n11), .B(any_edge), .Y(N24) );
  OAI21X1 U26 ( .B(n8), .C(n9), .A(n4), .Y(n14) );
  INVX1 U27 ( .A(dbcnt[11]), .Y(n4) );
  NAND3X1 U28 ( .A(dbcnt[8]), .B(dbcnt[10]), .C(dbcnt[9]), .Y(n9) );
  NOR42XL U29 ( .C(n8), .D(n15), .A(dbcnt[0]), .B(dbcnt[10]), .Y(n13) );
  NOR4XL U30 ( .A(dbcnt[9]), .B(dbcnt[8]), .C(dbcnt[2]), .D(dbcnt[1]), .Y(n15)
         );
  INVX1 U31 ( .A(n10), .Y(n8) );
  NAND32X1 U32 ( .B(dbcnt[4]), .C(dbcnt[3]), .A(n16), .Y(n10) );
  NOR3XL U33 ( .A(dbcnt[5]), .B(dbcnt[7]), .C(dbcnt[6]), .Y(n16) );
endmodule


module filter150us_a0_1_DW01_inc_0 ( A, SUM );
  input [11:0] A;
  output [11:0] SUM;

  wire   [11:2] carry;

  HAD1X1 U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .SO(SUM[10]) );
  HAD1X1 U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .SO(SUM[9]) );
  HAD1X1 U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .SO(SUM[8]) );
  HAD1X1 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .SO(SUM[7]) );
  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  XOR2X1 U1 ( .A(carry[11]), .B(A[11]), .Y(SUM[11]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_filter150us_a0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module ff_sync_0 ( i_org, o_dbc, o_chg, clk, rstz );
  input i_org, clk, rstz;
  output o_dbc, o_chg;
  wire   d_org_0_;

  DFFRQX1 d_org_reg_1_ ( .D(d_org_0_), .C(clk), .XR(rstz), .Q(o_dbc) );
  DFFRQX1 d_org_reg_0_ ( .D(i_org), .C(clk), .XR(rstz), .Q(d_org_0_) );
  XOR2X1 U3 ( .A(o_dbc), .B(d_org_0_), .Y(o_chg) );
endmodule


module ff_sync_1 ( i_org, o_dbc, o_chg, clk, rstz );
  input i_org, clk, rstz;
  output o_dbc, o_chg;
  wire   d_org_0_;

  DFFRQX1 d_org_reg_0_ ( .D(i_org), .C(clk), .XR(rstz), .Q(d_org_0_) );
  DFFRQX1 d_org_reg_1_ ( .D(d_org_0_), .C(clk), .XR(rstz), .Q(o_dbc) );
  XOR2X1 U3 ( .A(o_dbc), .B(d_org_0_), .Y(o_chg) );
endmodule


module ff_sync_2 ( i_org, o_dbc, o_chg, clk, rstz );
  input i_org, clk, rstz;
  output o_dbc, o_chg;
  wire   d_org_0_;

  DFFRQX1 d_org_reg_0_ ( .D(i_org), .C(clk), .XR(rstz), .Q(d_org_0_) );
  DFFRQX1 d_org_reg_1_ ( .D(d_org_0_), .C(clk), .XR(rstz), .Q(o_dbc) );
  XOR2X1 U3 ( .A(o_dbc), .B(d_org_0_), .Y(o_chg) );
endmodule


module dacmux_a0 ( clk, srstz, i_comp, r_comp_opt, r_wdat, r_adofs, r_isofs, 
        r_wr, dacv_wr, o_dacv, o_shrst, o_hold, o_dac1, o_daci_sel, o_dat, 
        r_dac_en, r_sar_en, o_dactl, o_cmpsta, x_daclsb, o_intr, o_smpl );
  input [2:0] r_comp_opt;
  input [7:0] r_wdat;
  output [7:0] r_adofs;
  output [7:0] r_isofs;
  input [10:0] r_wr;
  input [17:0] dacv_wr;
  output [143:0] o_dacv;
  output [9:0] o_dac1;
  output [17:0] o_daci_sel;
  output [17:0] o_dat;
  output [17:0] r_dac_en;
  output [17:0] r_sar_en;
  output [7:0] o_dactl;
  output [7:0] o_cmpsta;
  output [5:0] x_daclsb;
  output [4:0] o_smpl;
  input clk, srstz, i_comp;
  output o_shrst, o_hold, o_intr;
  wire   n534, n535, n536, n537, n538, n539, n540, n541, dacyc_done, updcmp,
         semi_start, auto_start, auto_sar, sacyc_done, sar_ini, sar_nxt,
         sampl_begn, sampl_done, ps_md4ch, ps_sample, updlsb, N859, tochg,
         N1239, N1240, N1241, N1242, N1243, N1244, N1245, N1246, N1247, N1250,
         N1251, N1252, N1253, N1254, N1255, N1256, N1257, N1258, N1261, N1262,
         N1263, N1264, N1265, N1266, N1267, N1268, N1269, N1272, N1273, N1274,
         N1275, N1276, N1277, N1278, N1279, N1280, N1283, N1284, N1285, N1286,
         N1287, N1288, N1289, N1290, N1291, N1294, N1295, N1296, N1297, N1298,
         N1299, N1300, N1301, N1302, N1305, N1306, N1307, N1308, N1309, N1310,
         N1311, N1312, N1313, N1316, N1317, N1318, N1319, N1320, N1321, N1322,
         N1323, N1324, N1327, N1328, N1329, N1330, N1331, N1332, N1333, N1334,
         N1335, N1338, N1339, N1340, N1341, N1342, N1343, N1344, N1345, N1346,
         N1349, N1350, N1351, N1352, N1353, N1354, N1355, N1356, N1357, N1360,
         N1361, N1362, N1363, N1364, N1365, N1366, N1367, N1368, N1371, N1372,
         N1373, N1374, N1375, N1376, N1377, N1378, N1379, N1382, N1383, N1384,
         N1385, N1386, N1387, N1388, N1389, N1390, N1393, N1394, N1395, N1396,
         N1397, N1398, N1399, N1400, N1401, N1404, N1405, N1406, N1407, N1408,
         N1409, N1410, N1411, N1412, N1415, N1416, N1417, N1418, N1419, N1420,
         N1421, N1422, N1423, N1426, N1427, N1428, N1429, N1430, N1431, N1432,
         N1433, N1434, n63, n98, n99, n101, n149, n150, n152, n159, n160, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n266,
         n267, n268, n270, n271, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n64, n65, n66, n67,
         n68, n69, n70, n72, n73, n74, n76, n78, n80, n82, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n100, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n151, n153, n154, n155, n156, n157, n158, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n265, n269, n272, n273, n274, n275, n276, n277, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533;
  wire   [1:0] syn_comp;
  wire   [4:0] cs_ptr;
  wire   [17:0] datcmp;
  wire   [4:0] ps_ptr;
  wire   [9:0] r_dac1v;
  wire   [9:0] r_rpt_v;
  wire   [17:0] app_dacis;
  wire   [17:0] pos_dacis;
  wire   [5:0] wdlsb;
  wire   [17:0] upd;
  wire   [7:0] wda;
  wire   [143:0] r_dacvs;
  wire   [7:0] setsta;
  wire   [7:0] clrsta;
  wire   [7:0] r_irq;

  glreg_00000012 u0_compi ( .clk(clk), .arstz(n163), .we(updcmp), .wdat(datcmp), .rdat(o_dat) );
  dac2sar_a0 u0_dac2sar ( .r_dac_t(o_dactl[3:2]), .r_dacyc(o_dactl[7]), 
        .r_sar10(n63), .sar_ini(sar_ini), .sar_nxt(sar_nxt), .semi_nxt(n99), 
        .auto_sar(auto_sar), .busy(o_dactl[0]), .stop(n19), .sync_i(
        syn_comp[1]), .sampl_begn(sampl_begn), .sampl_done(sampl_done), 
        .sh_rst(o_shrst), .dacyc_done(dacyc_done), .sacyc_done(sacyc_done), 
        .dac_v(r_dac1v), .rpt_v(r_rpt_v), .clk(clk), .srstz(srstz) );
  shmux_00000005_00000012_00000012 u0_shmux ( .ps_sample(ps_sample), 
        .ps_md4ch(ps_md4ch), .r_comp_swtch(r_comp_opt[2]), .r_semi(n101), 
        .r_loop(o_dactl[1]), .r_dac_en(r_dac_en), .wr_dacv(dacv_wr), .busy(
        o_dactl[0]), .sh_hold(o_hold), .stop(n19), .semi_start(semi_start), 
        .auto_start(auto_start), .mxcyc_done(n87), .sampl_begn(sampl_begn), 
        .sampl_done(sampl_done), .app_dacis(app_dacis), .pos_dacis(pos_dacis), 
        .cs_ptr(cs_ptr), .ps_ptr(ps_ptr), .clk(clk), .srstz(n171) );
  glreg_WIDTH7_1 u0_dactl ( .clk(clk), .arstz(n171), .we(n98), .wdat({
        r_wdat[7:6], n29, n26, r_wdat[3], n21, r_wdat[1]}), .rdat(o_dactl[7:1]) );
  glreg_a0_48 u0_dacen ( .clk(clk), .arstz(n141), .we(r_wr[1]), .wdat({
        r_wdat[7:6], n29, n26, r_wdat[3], n21, r_wdat[1], n118}), .rdat(
        r_dac_en[7:0]) );
  glreg_a0_47 u0_saren ( .clk(clk), .arstz(n142), .we(r_wr[2]), .wdat({
        r_wdat[7:6], n29, n26, r_wdat[3], n21, r_wdat[1], n119}), .rdat(
        r_sar_en[7:0]) );
  glreg_WIDTH6_2 u0_daclsb ( .clk(clk), .arstz(n172), .we(updlsb), .wdat(wdlsb), .rdat(x_daclsb) );
  glreg_a0_46 dacvs_0__u0 ( .clk(clk), .arstz(n143), .we(upd[0]), .wdat({n35, 
        n37, n38, n54, n40, n44, n62, n48}), .rdat(r_dacvs[7:0]) );
  glreg_a0_45 dacvs_1__u0 ( .clk(clk), .arstz(n157), .we(upd[1]), .wdat({n35, 
        n37, n39, n55, n41, n45, n85, n49}), .rdat(r_dacvs[15:8]) );
  glreg_a0_44 dacvs_2__u0 ( .clk(clk), .arstz(n144), .we(upd[2]), .wdat({n35, 
        n37, n39, n55, n41, n45, n85, n49}), .rdat(r_dacvs[23:16]) );
  glreg_a0_43 dacvs_3__u0 ( .clk(clk), .arstz(n145), .we(upd[3]), .wdat({
        wda[7:6], n38, n54, n40, n44, n85, n48}), .rdat(r_dacvs[31:24]) );
  glreg_a0_42 dacvs_4__u0 ( .clk(clk), .arstz(n146), .we(upd[4]), .wdat({n35, 
        n37, n39, n55, n41, n45, n85, n49}), .rdat(r_dacvs[39:32]) );
  glreg_a0_41 dacvs_5__u0 ( .clk(clk), .arstz(n147), .we(upd[5]), .wdat({
        wda[7:6], n39, n55, n41, n45, n62, n49}), .rdat(r_dacvs[47:40]) );
  glreg_a0_40 dacvs_6__u0 ( .clk(clk), .arstz(n148), .we(upd[6]), .wdat({
        wda[7:6], n39, n55, n41, n45, n62, n49}), .rdat(r_dacvs[55:48]) );
  glreg_a0_39 dacvs_7__u0 ( .clk(clk), .arstz(n151), .we(upd[7]), .wdat({
        wda[7:6], n39, n55, n41, n45, n62, n49}), .rdat(r_dacvs[63:56]) );
  glreg_a0_38 dacvs_8__u0 ( .clk(clk), .arstz(n153), .we(upd[8]), .wdat({
        wda[7:6], n39, n55, n41, n45, n85, n49}), .rdat(r_dacvs[71:64]) );
  glreg_a0_37 dacvs_9__u0 ( .clk(clk), .arstz(n154), .we(upd[9]), .wdat({
        wda[7:6], n39, n55, n41, n45, n62, n49}), .rdat(r_dacvs[79:72]) );
  glreg_a0_36 dacvs_10__u0 ( .clk(clk), .arstz(n155), .we(upd[10]), .wdat({
        wda[7:6], n38, n54, n40, n44, n62, n48}), .rdat(r_dacvs[87:80]) );
  glreg_a0_35 dacvs_11__u0 ( .clk(clk), .arstz(n156), .we(upd[11]), .wdat({
        wda[7:6], n39, n55, n41, n45, n85, n49}), .rdat(r_dacvs[95:88]) );
  glreg_a0_34 dacvs_12__u0 ( .clk(clk), .arstz(n158), .we(upd[12]), .wdat({
        wda[7:6], n38, n54, n40, n44, n85, n48}), .rdat(r_dacvs[103:96]) );
  glreg_a0_33 dacvs_13__u0 ( .clk(clk), .arstz(n161), .we(upd[13]), .wdat({n35, 
        n37, n38, n54, n40, n44, n62, n48}), .rdat(r_dacvs[111:104]) );
  glreg_a0_32 dacvs_14__u0 ( .clk(clk), .arstz(n162), .we(upd[14]), .wdat({n35, 
        n37, n38, n54, n40, n44, n85, n48}), .rdat(r_dacvs[119:112]) );
  glreg_a0_31 dacvs_15__u0 ( .clk(clk), .arstz(n163), .we(upd[15]), .wdat({n35, 
        n37, n38, n54, n40, n44, n62, n48}), .rdat(r_dacvs[127:120]) );
  glreg_a0_30 dacvs_16__u0 ( .clk(clk), .arstz(n164), .we(upd[16]), .wdat({n35, 
        n37, n38, n54, n40, n44, n62, n48}), .rdat(r_dacvs[135:128]) );
  glreg_a0_29 dacvs_17__u0 ( .clk(clk), .arstz(n165), .we(upd[17]), .wdat({n35, 
        n37, n38, n54, n40, n44, n85, n48}), .rdat(r_dacvs[143:136]) );
  glsta_a0_1 u0_cmpsta ( .clk(clk), .arstz(n166), .rst0(1'b0), .set2(setsta), 
        .clr1(clrsta), .rdat(o_cmpsta), .irq(r_irq) );
  glreg_a0_28 u0_adofs ( .clk(clk), .arstz(n167), .we(r_wr[5]), .wdat({
        r_wdat[7:6], n28, n25, r_wdat[3], n21, n23, n118}), .rdat({n534, n535, 
        n536, n537, n538, n539, n540, n541}) );
  glreg_a0_27 u0_isofs ( .clk(clk), .arstz(n168), .we(r_wr[6]), .wdat({
        r_wdat[7:6], n29, n26, r_wdat[3], n21, r_wdat[1], n119}), .rdat(
        r_isofs) );
  glreg_a0_26 u1_dacen ( .clk(clk), .arstz(n169), .we(r_wr[7]), .wdat({
        r_wdat[7:6], n29, n26, r_wdat[3], n21, r_wdat[1], n118}), .rdat(
        r_dac_en[15:8]) );
  glreg_a0_25 u1_saren ( .clk(clk), .arstz(n170), .we(r_wr[8]), .wdat({
        r_wdat[7:6], n29, n26, r_wdat[3], n21, r_wdat[1], n119}), .rdat(
        r_sar_en[15:8]) );
  glreg_WIDTH2_1 u2_dacen ( .clk(clk), .arstz(n172), .we(r_wr[9]), .wdat({
        r_wdat[1], n118}), .rdat(r_dac_en[17:16]) );
  glreg_WIDTH2_0 u2_saren ( .clk(clk), .arstz(n172), .we(r_wr[10]), .wdat({n23, 
        n119}), .rdat(r_sar_en[17:16]) );
  dacmux_a0_DW01_add_0 add_230_I18 ( .A({1'b0, r_dacvs[143:136]}), .B({n135, 
        n135, n535, n536, n537, n538, n539, n540, n31}), .CI(1'b0), .SUM({
        N1434, N1433, N1432, N1431, N1430, N1429, N1428, N1427, N1426}), .CO()
         );
  dacmux_a0_DW01_add_1 add_230_I17 ( .A({1'b0, r_dacvs[135:128]}), .B({n135, 
        n135, n535, n536, n537, n538, n539, n540, n33}), .CI(1'b0), .SUM({
        N1423, N1422, N1421, N1420, N1419, N1418, N1417, N1416, N1415}), .CO()
         );
  dacmux_a0_DW01_add_2 add_230_I16 ( .A({1'b0, r_dacvs[127:120]}), .B({n135, 
        n135, r_adofs[6:1], n33}), .CI(1'b0), .SUM({N1412, N1411, N1410, N1409, 
        N1408, N1407, N1406, N1405, N1404}), .CO() );
  dacmux_a0_DW01_add_3 add_230_I15 ( .A({1'b0, r_dacvs[119:112]}), .B({n135, 
        n135, r_adofs[6:1], n31}), .CI(1'b0), .SUM({N1401, N1400, N1399, N1398, 
        N1397, N1396, N1395, N1394, N1393}), .CO() );
  dacmux_a0_DW01_add_4 add_230_I14 ( .A({1'b0, r_dacvs[111:104]}), .B({n135, 
        n135, r_adofs[6:1], n541}), .CI(1'b0), .SUM({N1390, N1389, N1388, 
        N1387, N1386, N1385, N1384, N1383, N1382}), .CO() );
  dacmux_a0_DW01_add_5 add_230_I13 ( .A({1'b0, r_dacvs[103:96]}), .B({n136, 
        n136, n535, n536, n537, n538, n539, n540, r_adofs[0]}), .CI(1'b0), 
        .SUM({N1379, N1378, N1377, N1376, N1375, N1374, N1373, N1372, N1371}), 
        .CO() );
  dacmux_a0_DW01_add_6 add_230_I12 ( .A({1'b0, r_dacvs[95:88]}), .B({n136, 
        n136, n535, n536, n537, n538, n539, n540, n541}), .CI(1'b0), .SUM({
        N1368, N1367, N1366, N1365, N1364, N1363, N1362, N1361, N1360}), .CO()
         );
  dacmux_a0_DW01_add_7 add_230_I11 ( .A({1'b0, r_dacvs[87:80]}), .B({n136, 
        n136, n535, n536, n537, n538, n539, n540, n33}), .CI(1'b0), .SUM({
        N1357, N1356, N1355, N1354, N1353, N1352, N1351, N1350, N1349}), .CO()
         );
  dacmux_a0_DW01_add_8 add_230_I10 ( .A({1'b0, r_dacvs[79:72]}), .B({n136, 
        n136, r_adofs[6:1], n31}), .CI(1'b0), .SUM({N1346, N1345, N1344, N1343, 
        N1342, N1341, N1340, N1339, N1338}), .CO() );
  dacmux_a0_DW01_add_9 add_230_I9 ( .A({1'b0, r_dacvs[71:64]}), .B({n136, n137, 
        n535, n536, n537, n538, n539, n540, r_adofs[0]}), .CI(1'b0), .SUM({
        N1335, N1334, N1333, N1332, N1331, N1330, N1329, N1328, N1327}), .CO()
         );
  dacmux_a0_DW01_add_10 add_230_I8 ( .A({1'b0, r_dacvs[63:56]}), .B({n137, 
        n137, r_adofs[6:0]}), .CI(1'b0), .SUM({N1324, N1323, N1322, N1321, 
        N1320, N1319, N1318, N1317, N1316}), .CO() );
  dacmux_a0_DW01_add_11 add_230_I7 ( .A({1'b0, r_dacvs[55:48]}), .B({n137, 
        n137, n535, n536, n537, n538, n539, n540, n33}), .CI(1'b0), .SUM({
        N1313, N1312, N1311, N1310, N1309, N1308, N1307, N1306, N1305}), .CO()
         );
  dacmux_a0_DW01_add_12 add_230_I6 ( .A({1'b0, r_dacvs[47:40]}), .B({n137, 
        n137, r_adofs[6:1], n33}), .CI(1'b0), .SUM({N1302, N1301, N1300, N1299, 
        N1298, N1297, N1296, N1295, N1294}), .CO() );
  dacmux_a0_DW01_add_13 add_230_I5 ( .A({1'b0, r_dacvs[39:32]}), .B({n137, 
        n137, r_adofs[6:1], n31}), .CI(1'b0), .SUM({N1291, N1290, N1289, N1288, 
        N1287, N1286, N1285, N1284, N1283}), .CO() );
  dacmux_a0_DW01_add_14 add_230_I4 ( .A({1'b0, r_dacvs[31:24]}), .B({n137, 
        r_adofs[7], n535, n536, n537, n538, n539, n540, r_adofs[0]}), .CI(1'b0), .SUM({N1280, N1279, N1278, N1277, N1276, N1275, N1274, N1273, N1272}), .CO()
         );
  dacmux_a0_DW01_add_15 add_230_I3 ( .A({1'b0, r_dacvs[23:16]}), .B({
        r_isofs[7], r_isofs}), .CI(1'b0), .SUM({N1269, N1268, N1267, N1266, 
        N1265, N1264, N1263, N1262, N1261}), .CO() );
  dacmux_a0_DW01_add_16 add_230_I2 ( .A({1'b0, r_dacvs[15:8]}), .B({r_adofs[7], 
        r_adofs[7:1], n31}), .CI(1'b0), .SUM({N1258, N1257, N1256, N1255, 
        N1254, N1253, N1252, N1251, N1250}), .CO() );
  dacmux_a0_DW01_add_17 add_230 ( .A({1'b0, r_dacvs[7:0]}), .B({r_adofs[7], 
        n136, n535, n536, n537, n538, n539, n540, n541}), .CI(1'b0), .SUM({
        N1247, N1246, N1245, N1244, N1243, N1242, N1241, N1240, N1239}), .CO()
         );
  DFFQX1 syn_comp_reg_1_ ( .D(syn_comp[0]), .C(clk), .Q(syn_comp[1]) );
  DFFQX1 syn_comp_reg_0_ ( .D(i_comp), .C(clk), .Q(syn_comp[0]) );
  NAND21X1 U3 ( .B(ps_ptr[4]), .A(n409), .Y(n385) );
  NOR21XL U4 ( .B(r_dac_en[16]), .A(n382), .Y(n392) );
  MUX2IX1 U5 ( .D0(n390), .D1(n389), .S(ps_ptr[3]), .Y(n391) );
  MUX2IX1 U6 ( .D0(n415), .D1(n414), .S(ps_ptr[0]), .Y(n416) );
  AO21X1 U7 ( .B(N1253), .C(n459), .A(n458), .Y(o_dacv[11]) );
  INVX1 U8 ( .A(n384), .Y(n409) );
  INVX1 U9 ( .A(n388), .Y(n406) );
  AO2222XL U10 ( .A(r_dac_en[8]), .B(n409), .C(r_dac_en[10]), .D(n408), .E(
        r_dac_en[12]), .F(n407), .G(r_dac_en[14]), .H(n406), .Y(n389) );
  INVX2 U11 ( .A(n399), .Y(auto_start) );
  NAND21X1 U12 ( .B(n419), .A(n418), .Y(n420) );
  NOR21XL U13 ( .B(n417), .A(n416), .Y(n418) );
  INVX1 U14 ( .A(r_wdat[0]), .Y(n86) );
  AND2X1 U15 ( .A(n86), .B(r_wr[0]), .Y(n19) );
  INVX1 U16 ( .A(r_wdat[2]), .Y(n20) );
  INVX1 U17 ( .A(n20), .Y(n21) );
  INVX1 U18 ( .A(r_wdat[1]), .Y(n22) );
  INVX1 U19 ( .A(n22), .Y(n23) );
  INVX1 U20 ( .A(r_wdat[4]), .Y(n24) );
  INVX1 U21 ( .A(n24), .Y(n25) );
  INVX1 U22 ( .A(n24), .Y(n26) );
  INVX1 U23 ( .A(r_wdat[5]), .Y(n27) );
  INVX1 U42 ( .A(n27), .Y(n28) );
  INVX1 U43 ( .A(n27), .Y(n29) );
  INVX1 U44 ( .A(n541), .Y(n30) );
  INVX1 U45 ( .A(n30), .Y(n31) );
  INVX1 U46 ( .A(n30), .Y(r_adofs[0]) );
  INVX1 U47 ( .A(n30), .Y(n33) );
  INVX1 U48 ( .A(wda[7]), .Y(n34) );
  INVX1 U49 ( .A(n34), .Y(n35) );
  INVX1 U50 ( .A(wda[6]), .Y(n36) );
  INVX1 U51 ( .A(n36), .Y(n37) );
  BUFX3 U52 ( .A(n424), .Y(wda[5]) );
  INVX1 U53 ( .A(wda[5]), .Y(n38) );
  INVX1 U54 ( .A(wda[5]), .Y(n39) );
  BUFX3 U55 ( .A(n427), .Y(wda[3]) );
  INVX1 U56 ( .A(wda[3]), .Y(n40) );
  INVX1 U57 ( .A(wda[3]), .Y(n41) );
  NAND2X1 U58 ( .A(n378), .B(n199), .Y(n298) );
  INVX1 U59 ( .A(n298), .Y(n42) );
  INVX1 U60 ( .A(n298), .Y(n43) );
  BUFX3 U61 ( .A(n428), .Y(wda[2]) );
  INVX1 U62 ( .A(wda[2]), .Y(n44) );
  INVX1 U63 ( .A(wda[2]), .Y(n45) );
  NAND2X1 U64 ( .A(n378), .B(n375), .Y(n294) );
  INVX1 U65 ( .A(n294), .Y(n46) );
  INVX1 U66 ( .A(n294), .Y(n47) );
  BUFX3 U67 ( .A(n430), .Y(wda[0]) );
  INVX1 U68 ( .A(wda[0]), .Y(n48) );
  INVX1 U69 ( .A(wda[0]), .Y(n49) );
  NAND2X1 U70 ( .A(n374), .B(n199), .Y(n296) );
  INVX1 U71 ( .A(n296), .Y(n50) );
  INVX1 U72 ( .A(n296), .Y(n51) );
  NAND2X1 U73 ( .A(n377), .B(n375), .Y(n291) );
  INVX1 U74 ( .A(n291), .Y(n52) );
  INVX1 U75 ( .A(n291), .Y(n53) );
  BUFX3 U76 ( .A(n425), .Y(wda[4]) );
  INVX1 U77 ( .A(wda[4]), .Y(n54) );
  INVX1 U78 ( .A(wda[4]), .Y(n55) );
  INVX1 U79 ( .A(n379), .Y(n56) );
  NAND2X1 U80 ( .A(n377), .B(n199), .Y(n297) );
  INVX1 U81 ( .A(n297), .Y(n57) );
  INVX1 U82 ( .A(n297), .Y(n58) );
  NAND2X1 U83 ( .A(n375), .B(n376), .Y(n292) );
  INVX1 U84 ( .A(n292), .Y(n59) );
  INVX1 U85 ( .A(n292), .Y(n60) );
  INVX1 U86 ( .A(n85), .Y(n61) );
  INVX1 U87 ( .A(n61), .Y(n62) );
  NAND21X2 U88 ( .B(n421), .A(n420), .Y(sar_ini) );
  NAND2X1 U89 ( .A(n376), .B(n199), .Y(n295) );
  INVX1 U90 ( .A(n295), .Y(n64) );
  INVX1 U91 ( .A(n295), .Y(n65) );
  NAND2X1 U92 ( .A(n374), .B(n375), .Y(n293) );
  INVX1 U93 ( .A(n293), .Y(n66) );
  INVX1 U94 ( .A(n293), .Y(n67) );
  BUFX3 U95 ( .A(n299), .Y(n68) );
  INVX1 U96 ( .A(r_comp_opt[0]), .Y(n120) );
  INVX1 U97 ( .A(n120), .Y(n69) );
  INVX1 U98 ( .A(n535), .Y(n70) );
  INVX1 U99 ( .A(n70), .Y(r_adofs[6]) );
  NOR2X1 U100 ( .A(o_dactl[0]), .B(semi_start), .Y(n453) );
  INVX1 U101 ( .A(n453), .Y(n72) );
  INVX1 U102 ( .A(n453), .Y(n73) );
  INVX1 U103 ( .A(n537), .Y(n74) );
  INVX1 U104 ( .A(n74), .Y(r_adofs[4]) );
  INVX1 U105 ( .A(n536), .Y(n76) );
  INVX1 U106 ( .A(n76), .Y(r_adofs[5]) );
  INVX1 U107 ( .A(n539), .Y(n78) );
  INVX1 U108 ( .A(n78), .Y(r_adofs[2]) );
  INVX1 U109 ( .A(n540), .Y(n80) );
  INVX1 U110 ( .A(n80), .Y(r_adofs[1]) );
  INVX1 U111 ( .A(n538), .Y(n82) );
  INVX1 U112 ( .A(n82), .Y(r_adofs[3]) );
  AO2222X1 U113 ( .A(n409), .B(r_sar_en[9]), .C(n408), .D(r_sar_en[11]), .E(
        n407), .F(r_sar_en[13]), .G(n406), .H(r_sar_en[15]), .Y(n410) );
  INVXL U114 ( .A(dacv_wr[15]), .Y(n433) );
  NAND21XL U115 ( .B(n387), .A(ps_ptr[2]), .Y(n388) );
  NAND21XL U116 ( .B(n421), .A(n381), .Y(semi_start) );
  INVX2 U117 ( .A(n386), .Y(n407) );
  AND2XL U118 ( .A(n23), .B(r_wr[4]), .Y(clrsta[1]) );
  AND4X1 U119 ( .A(n196), .B(n195), .C(n194), .D(n84), .Y(n197) );
  AOI22XL U120 ( .A(dacv_wr[17]), .B(r_sar_en[17]), .C(dacv_wr[16]), .D(
        r_sar_en[16]), .Y(n84) );
  MUX2BXL U121 ( .D0(r_rpt_v[3]), .D1(n22), .S(n121), .Y(n85) );
  INVX1 U122 ( .A(dacv_wr[4]), .Y(n447) );
  INVX1 U123 ( .A(dacv_wr[5]), .Y(n445) );
  INVX1 U124 ( .A(n125), .Y(n117) );
  INVX1 U125 ( .A(n125), .Y(n116) );
  INVX1 U126 ( .A(n173), .Y(n172) );
  INVX1 U127 ( .A(n173), .Y(n166) );
  INVX1 U128 ( .A(n173), .Y(n165) );
  INVX1 U129 ( .A(n174), .Y(n164) );
  INVX1 U130 ( .A(n175), .Y(n163) );
  INVX1 U131 ( .A(n175), .Y(n162) );
  INVX1 U132 ( .A(n174), .Y(n161) );
  INVX1 U133 ( .A(n173), .Y(n158) );
  INVX1 U134 ( .A(n174), .Y(n156) );
  INVX1 U135 ( .A(n174), .Y(n155) );
  INVX1 U136 ( .A(n175), .Y(n154) );
  INVX1 U137 ( .A(n173), .Y(n153) );
  INVX1 U138 ( .A(n174), .Y(n151) );
  INVX1 U139 ( .A(n175), .Y(n148) );
  INVX1 U140 ( .A(n174), .Y(n147) );
  INVX1 U141 ( .A(n174), .Y(n146) );
  INVX1 U142 ( .A(n175), .Y(n145) );
  INVX1 U143 ( .A(n175), .Y(n144) );
  INVX1 U144 ( .A(n175), .Y(n157) );
  INVX1 U145 ( .A(n175), .Y(n143) );
  INVX1 U146 ( .A(n174), .Y(n170) );
  INVX1 U147 ( .A(n174), .Y(n169) );
  INVX1 U148 ( .A(n174), .Y(n168) );
  INVX1 U149 ( .A(n173), .Y(n167) );
  INVX1 U150 ( .A(n175), .Y(n142) );
  INVX1 U151 ( .A(n173), .Y(n171) );
  INVX1 U152 ( .A(dacv_wr[13]), .Y(n435) );
  INVX1 U153 ( .A(dacv_wr[6]), .Y(n444) );
  INVX1 U154 ( .A(srstz), .Y(n173) );
  INVX1 U155 ( .A(r_wr[3]), .Y(n491) );
  INVX1 U156 ( .A(r_wr[4]), .Y(n490) );
  INVX1 U157 ( .A(n492), .Y(n121) );
  INVX1 U158 ( .A(n492), .Y(n122) );
  NOR2X1 U159 ( .A(n126), .B(n128), .Y(n378) );
  INVX1 U160 ( .A(n492), .Y(n123) );
  NAND2X1 U161 ( .A(n124), .B(n126), .Y(n532) );
  NAND21X1 U162 ( .B(n126), .A(n124), .Y(n450) );
  NAND21X1 U163 ( .B(n124), .A(n126), .Y(n449) );
  NAND21X1 U164 ( .B(n451), .A(n446), .Y(n498) );
  NAND21X1 U165 ( .B(n450), .A(n446), .Y(n511) );
  NAND21X1 U166 ( .B(n451), .A(n441), .Y(n499) );
  NAND21X1 U167 ( .B(n450), .A(n441), .Y(n512) );
  NAND21X1 U168 ( .B(n451), .A(n431), .Y(n497) );
  NAND21X1 U169 ( .B(n450), .A(n431), .Y(n509) );
  NAND21X1 U170 ( .B(n449), .A(n446), .Y(n503) );
  NAND21X1 U171 ( .B(n448), .A(n446), .Y(n507) );
  NAND21X1 U172 ( .B(n449), .A(n441), .Y(n500) );
  NAND21X1 U173 ( .B(n448), .A(n441), .Y(n504) );
  OR2X1 U174 ( .A(n452), .B(n451), .Y(n495) );
  OR2X1 U175 ( .A(n452), .B(n450), .Y(n510) );
  OR2X1 U176 ( .A(n452), .B(n449), .Y(n502) );
  OR2X1 U177 ( .A(n452), .B(n448), .Y(n506) );
  INVX1 U178 ( .A(n175), .Y(n141) );
  INVX1 U179 ( .A(srstz), .Y(n175) );
  INVX1 U180 ( .A(srstz), .Y(n174) );
  NAND21X1 U181 ( .B(ps_ptr[2]), .A(n387), .Y(n384) );
  INVX1 U182 ( .A(n381), .Y(n99) );
  NOR2X1 U183 ( .A(n479), .B(n490), .Y(clrsta[6]) );
  NOR2X1 U184 ( .A(n478), .B(n490), .Y(clrsta[7]) );
  INVX1 U185 ( .A(n125), .Y(n124) );
  NOR2X1 U186 ( .A(n533), .B(n529), .Y(setsta[4]) );
  NOR2X1 U187 ( .A(n533), .B(n530), .Y(setsta[5]) );
  NOR2X1 U188 ( .A(n533), .B(n531), .Y(setsta[6]) );
  INVX1 U189 ( .A(n130), .Y(n115) );
  NOR2X1 U190 ( .A(n533), .B(n532), .Y(setsta[7]) );
  INVX1 U191 ( .A(n127), .Y(n126) );
  NOR2X1 U192 ( .A(n56), .B(n124), .Y(n285) );
  INVX1 U193 ( .A(n129), .Y(n128) );
  NOR2X1 U194 ( .A(n129), .B(n126), .Y(n374) );
  NOR2X1 U195 ( .A(n127), .B(n128), .Y(n376) );
  INVX1 U196 ( .A(n130), .Y(n114) );
  NOR2X1 U197 ( .A(n127), .B(n129), .Y(n377) );
  NAND2X1 U198 ( .A(n126), .B(n125), .Y(n531) );
  NAND2X1 U199 ( .A(n124), .B(n127), .Y(n530) );
  NAND21X1 U200 ( .B(n124), .A(n127), .Y(n451) );
  NAND21X1 U201 ( .B(n127), .A(n124), .Y(n448) );
  NAND32X1 U202 ( .B(n131), .C(n128), .A(n130), .Y(n452) );
  NAND21X1 U203 ( .B(n451), .A(n88), .Y(n496) );
  NAND21X1 U204 ( .B(n450), .A(n88), .Y(n508) );
  NAND21X1 U205 ( .B(n449), .A(n88), .Y(n501) );
  NAND21X1 U206 ( .B(n448), .A(n88), .Y(n505) );
  INVX1 U207 ( .A(n443), .Y(n446) );
  NAND32X1 U208 ( .B(n131), .C(n129), .A(n130), .Y(n443) );
  INVX1 U209 ( .A(n437), .Y(n441) );
  NAND32X1 U210 ( .B(n128), .C(n130), .A(n132), .Y(n437) );
  INVX1 U211 ( .A(n422), .Y(n431) );
  NAND32X1 U212 ( .B(n128), .C(n132), .A(n130), .Y(n422) );
  INVX1 U213 ( .A(ps_ptr[1]), .Y(n387) );
  NAND21XL U214 ( .B(ps_ptr[1]), .A(ps_ptr[2]), .Y(n386) );
  INVX1 U215 ( .A(n276), .Y(n421) );
  INVX1 U216 ( .A(r_wdat[3]), .Y(n426) );
  INVX1 U217 ( .A(N1313), .Y(n474) );
  INVX1 U218 ( .A(N1324), .Y(n477) );
  INVX1 U219 ( .A(N1258), .Y(n459) );
  INVX1 U220 ( .A(N1280), .Y(n465) );
  INVX1 U221 ( .A(n472), .Y(n473) );
  NAND21X1 U222 ( .B(r_adofs[7]), .A(N1313), .Y(n472) );
  INVX1 U223 ( .A(n475), .Y(n476) );
  NAND21X1 U224 ( .B(r_adofs[7]), .A(N1324), .Y(n475) );
  INVX1 U225 ( .A(n457), .Y(n458) );
  NAND21X1 U226 ( .B(r_adofs[7]), .A(N1258), .Y(n457) );
  INVX1 U227 ( .A(n454), .Y(n455) );
  NAND21X1 U228 ( .B(r_adofs[7]), .A(N1247), .Y(n454) );
  INVX1 U229 ( .A(n463), .Y(n464) );
  NAND21X1 U230 ( .B(r_adofs[7]), .A(N1280), .Y(n463) );
  OAI22X1 U231 ( .A(n432), .B(n72), .C(n497), .D(n123), .Y(upd[16]) );
  INVXL U232 ( .A(dacv_wr[16]), .Y(n432) );
  OAI22X1 U233 ( .A(n433), .B(n72), .C(n505), .D(n123), .Y(upd[15]) );
  OAI22X1 U234 ( .A(n434), .B(n72), .C(n501), .D(n123), .Y(upd[14]) );
  OAI22X1 U235 ( .A(n435), .B(n72), .C(n508), .D(n123), .Y(upd[13]) );
  OAI22X1 U236 ( .A(n436), .B(n72), .C(n496), .D(n123), .Y(upd[12]) );
  OAI22X1 U237 ( .A(n438), .B(n72), .C(n504), .D(n122), .Y(upd[11]) );
  INVXL U238 ( .A(dacv_wr[11]), .Y(n438) );
  OAI22X1 U239 ( .A(n439), .B(n72), .C(n500), .D(n122), .Y(upd[10]) );
  OAI22X1 U240 ( .A(n440), .B(n72), .C(n512), .D(n122), .Y(upd[9]) );
  INVXL U241 ( .A(dacv_wr[9]), .Y(n440) );
  OAI22X1 U242 ( .A(n442), .B(n72), .C(n499), .D(n122), .Y(upd[8]) );
  INVXL U243 ( .A(dacv_wr[8]), .Y(n442) );
  OAI22AX1 U244 ( .D(dacv_wr[7]), .C(n73), .A(n507), .B(n122), .Y(upd[7]) );
  OAI22X1 U245 ( .A(n444), .B(n73), .C(n503), .D(n122), .Y(upd[6]) );
  OAI22X1 U246 ( .A(n445), .B(n73), .C(n511), .D(n122), .Y(upd[5]) );
  OAI22X1 U247 ( .A(n447), .B(n73), .C(n498), .D(n122), .Y(upd[4]) );
  OAI22AX1 U248 ( .D(dacv_wr[3]), .C(n73), .A(n506), .B(n122), .Y(upd[3]) );
  OAI22AX1 U249 ( .D(dacv_wr[1]), .C(n73), .A(n510), .B(n122), .Y(upd[1]) );
  OAI22X1 U250 ( .A(n423), .B(n73), .C(n509), .D(n121), .Y(upd[17]) );
  INVXL U251 ( .A(dacv_wr[17]), .Y(n423) );
  OAI22AX1 U252 ( .D(dacv_wr[2]), .C(n73), .A(n502), .B(n121), .Y(upd[2]) );
  OAI22AX1 U253 ( .D(dacv_wr[0]), .C(n73), .A(n495), .B(n121), .Y(upd[0]) );
  INVX1 U254 ( .A(N1379), .Y(n484) );
  INVX1 U255 ( .A(N1434), .Y(n489) );
  INVX1 U256 ( .A(N1423), .Y(n488) );
  INVX1 U257 ( .A(N1346), .Y(n481) );
  INVX1 U258 ( .A(N1335), .Y(n480) );
  INVX1 U259 ( .A(N1412), .Y(n487) );
  INVX1 U260 ( .A(N1368), .Y(n483) );
  INVX1 U261 ( .A(N1357), .Y(n482) );
  INVX1 U262 ( .A(N1401), .Y(n486) );
  INVX1 U263 ( .A(N1390), .Y(n485) );
  INVX1 U264 ( .A(N1291), .Y(n468) );
  INVX1 U265 ( .A(N1302), .Y(n471) );
  INVX1 U266 ( .A(N1247), .Y(n456) );
  INVX1 U267 ( .A(n466), .Y(n467) );
  NAND21X1 U268 ( .B(n534), .A(N1291), .Y(n466) );
  INVX1 U269 ( .A(n469), .Y(n470) );
  NAND21X1 U270 ( .B(n534), .A(N1302), .Y(n469) );
  INVX1 U271 ( .A(r_wdat[6]), .Y(n479) );
  AND2X1 U272 ( .A(n29), .B(r_wr[4]), .Y(clrsta[5]) );
  AND2X1 U273 ( .A(n21), .B(r_wr[4]), .Y(clrsta[2]) );
  AND2X1 U274 ( .A(n26), .B(r_wr[4]), .Y(clrsta[4]) );
  AND2X1 U275 ( .A(r_wdat[3]), .B(r_wr[4]), .Y(clrsta[3]) );
  INVX1 U276 ( .A(r_wdat[7]), .Y(n478) );
  OA21X1 U277 ( .B(n243), .C(n520), .A(n244), .Y(n239) );
  AND2X1 U278 ( .A(n231), .B(n237), .Y(n238) );
  NOR2X1 U279 ( .A(n239), .B(n241), .Y(n242) );
  MUX2AXL U280 ( .D0(n494), .D1(sacyc_done), .S(auto_sar), .Y(n87) );
  INVX1 U281 ( .A(cs_ptr[0]), .Y(n125) );
  OR3XL U282 ( .A(n528), .B(cs_ptr[3]), .C(n131), .Y(n533) );
  NOR2X1 U283 ( .A(n529), .B(n527), .Y(setsta[0]) );
  NOR2X1 U284 ( .A(n531), .B(n527), .Y(setsta[2]) );
  NOR2X1 U285 ( .A(n530), .B(n527), .Y(setsta[1]) );
  NOR2X1 U286 ( .A(n532), .B(n527), .Y(setsta[3]) );
  INVX1 U287 ( .A(cs_ptr[1]), .Y(n127) );
  AND2X1 U288 ( .A(n124), .B(n379), .Y(n283) );
  INVX1 U289 ( .A(n132), .Y(n131) );
  INVX1 U290 ( .A(cs_ptr[4]), .Y(n132) );
  NOR2X1 U291 ( .A(cs_ptr[3]), .B(n131), .Y(n199) );
  INVX1 U292 ( .A(n379), .Y(n493) );
  INVX1 U293 ( .A(cs_ptr[2]), .Y(n129) );
  INVX1 U294 ( .A(dacyc_done), .Y(n494) );
  NOR32XL U295 ( .B(n378), .C(n131), .A(cs_ptr[3]), .Y(n299) );
  NOR21XL U296 ( .B(cs_ptr[3]), .A(n131), .Y(n375) );
  AO21X1 U297 ( .B(n101), .C(dacyc_done), .A(sacyc_done), .Y(n492) );
  NAND21X1 U298 ( .B(cs_ptr[0]), .A(n127), .Y(n529) );
  NOR31X1 U299 ( .C(cs_ptr[2]), .A(n130), .B(cs_ptr[4]), .Y(n88) );
  INVX1 U300 ( .A(cs_ptr[3]), .Y(n130) );
  AO21X1 U301 ( .B(N1240), .C(n456), .A(n455), .Y(o_dacv[1]) );
  AO21X1 U302 ( .B(N1265), .C(n462), .A(n461), .Y(o_dacv[20]) );
  AO21X1 U303 ( .B(N1266), .C(n462), .A(n461), .Y(o_dacv[21]) );
  AO21X1 U304 ( .B(N1267), .C(n462), .A(n461), .Y(o_dacv[22]) );
  AO21X1 U305 ( .B(N1244), .C(n456), .A(n455), .Y(o_dacv[5]) );
  AO21X1 U306 ( .B(N1245), .C(n456), .A(n455), .Y(o_dacv[6]) );
  AO21X1 U307 ( .B(N1287), .C(n468), .A(n467), .Y(o_dacv[36]) );
  AO21X1 U308 ( .B(N1284), .C(n468), .A(n467), .Y(o_dacv[33]) );
  AO21X1 U309 ( .B(N1296), .C(n471), .A(n470), .Y(o_dacv[42]) );
  AO21X1 U310 ( .B(N1298), .C(n471), .A(n470), .Y(o_dacv[44]) );
  AO21X1 U311 ( .B(N1295), .C(n471), .A(n470), .Y(o_dacv[41]) );
  AO21X1 U312 ( .B(N1297), .C(n471), .A(n470), .Y(o_dacv[43]) );
  AO21X1 U313 ( .B(N1274), .C(n465), .A(n464), .Y(o_dacv[26]) );
  AO21X1 U314 ( .B(N1276), .C(n465), .A(n464), .Y(o_dacv[28]) );
  AO21X1 U315 ( .B(N1273), .C(n465), .A(n464), .Y(o_dacv[25]) );
  AO21X1 U316 ( .B(N1275), .C(n465), .A(n464), .Y(o_dacv[27]) );
  AO21X1 U317 ( .B(N1290), .C(n468), .A(n467), .Y(o_dacv[39]) );
  INVX1 U318 ( .A(o_dactl[0]), .Y(n186) );
  NOR32XL U319 ( .B(n275), .C(n274), .A(n273), .Y(n277) );
  NOR32XL U320 ( .B(n272), .C(n269), .A(n265), .Y(n273) );
  AO21X1 U321 ( .B(N1309), .C(n474), .A(n473), .Y(o_dacv[52]) );
  AO21X1 U322 ( .B(N1320), .C(n477), .A(n476), .Y(o_dacv[60]) );
  AO21X1 U323 ( .B(N1242), .C(n456), .A(n455), .Y(o_dacv[3]) );
  AO21X1 U324 ( .B(N1243), .C(n456), .A(n455), .Y(o_dacv[4]) );
  AO21X1 U325 ( .B(N1321), .C(n477), .A(n476), .Y(o_dacv[61]) );
  AO21X1 U326 ( .B(N1306), .C(n474), .A(n473), .Y(o_dacv[49]) );
  AO21X1 U327 ( .B(N1241), .C(n456), .A(n455), .Y(o_dacv[2]) );
  AO21X1 U328 ( .B(N1246), .C(n456), .A(n455), .Y(o_dacv[7]) );
  AO21X1 U329 ( .B(N1286), .C(n468), .A(n467), .Y(o_dacv[35]) );
  AO21X1 U330 ( .B(N1299), .C(n471), .A(n470), .Y(o_dacv[45]) );
  AO21X1 U331 ( .B(N1288), .C(n468), .A(n467), .Y(o_dacv[37]) );
  AO21X1 U332 ( .B(N1289), .C(n468), .A(n467), .Y(o_dacv[38]) );
  AO21X1 U333 ( .B(N1300), .C(n471), .A(n470), .Y(o_dacv[46]) );
  AO21X1 U334 ( .B(N1285), .C(n468), .A(n467), .Y(o_dacv[34]) );
  AO21X1 U335 ( .B(N1322), .C(n477), .A(n476), .Y(o_dacv[62]) );
  AO21X1 U336 ( .B(N1301), .C(n471), .A(n470), .Y(o_dacv[47]) );
  NAND2X1 U337 ( .A(N1379), .B(n139), .Y(n266) );
  NAND2X1 U338 ( .A(N1423), .B(n140), .Y(n279) );
  NAND2X1 U339 ( .A(N1412), .B(n139), .Y(n280) );
  NAND2X1 U340 ( .A(N1401), .B(n140), .Y(n281) );
  NAND2X1 U341 ( .A(N1390), .B(n139), .Y(n282) );
  OAI21BBX1 U342 ( .A(N1367), .B(n483), .C(n267), .Y(o_dacv[95]) );
  OAI21BBX1 U343 ( .A(N1356), .B(n482), .C(n268), .Y(o_dacv[87]) );
  OAI21BBX1 U344 ( .A(N1400), .B(n486), .C(n281), .Y(o_dacv[119]) );
  OAI21BBX1 U345 ( .A(N1378), .B(n484), .C(n266), .Y(o_dacv[103]) );
  OAI21BBX1 U346 ( .A(N1389), .B(n485), .C(n282), .Y(o_dacv[111]) );
  OAI21BBX1 U347 ( .A(N1365), .B(n483), .C(n267), .Y(o_dacv[93]) );
  OAI21BBX1 U348 ( .A(N1354), .B(n482), .C(n268), .Y(o_dacv[85]) );
  OAI21BBX1 U349 ( .A(N1398), .B(n486), .C(n281), .Y(o_dacv[117]) );
  OAI21BBX1 U350 ( .A(N1376), .B(n484), .C(n266), .Y(o_dacv[101]) );
  OAI21BBX1 U351 ( .A(N1387), .B(n485), .C(n282), .Y(o_dacv[109]) );
  OAI21BBX1 U352 ( .A(N1366), .B(n483), .C(n267), .Y(o_dacv[94]) );
  OAI21BBX1 U353 ( .A(N1355), .B(n482), .C(n268), .Y(o_dacv[86]) );
  OAI21BBX1 U354 ( .A(N1399), .B(n486), .C(n281), .Y(o_dacv[118]) );
  OAI21BBX1 U355 ( .A(N1377), .B(n484), .C(n266), .Y(o_dacv[102]) );
  OAI21BBX1 U356 ( .A(N1388), .B(n485), .C(n282), .Y(o_dacv[110]) );
  OAI21BBX1 U357 ( .A(N1364), .B(n483), .C(n267), .Y(o_dacv[92]) );
  OAI21BBX1 U358 ( .A(N1353), .B(n482), .C(n268), .Y(o_dacv[84]) );
  OAI21BBX1 U359 ( .A(N1397), .B(n486), .C(n281), .Y(o_dacv[116]) );
  OAI21BBX1 U360 ( .A(N1375), .B(n484), .C(n266), .Y(o_dacv[100]) );
  OAI21BBX1 U361 ( .A(N1363), .B(n483), .C(n267), .Y(o_dacv[91]) );
  OAI21BBX1 U362 ( .A(N1352), .B(n482), .C(n268), .Y(o_dacv[83]) );
  OAI21BBX1 U363 ( .A(N1396), .B(n486), .C(n281), .Y(o_dacv[115]) );
  OAI21BBX1 U364 ( .A(N1374), .B(n484), .C(n266), .Y(o_dacv[99]) );
  OAI21BBX1 U365 ( .A(N1385), .B(n485), .C(n282), .Y(o_dacv[107]) );
  OAI21BBX1 U366 ( .A(N1362), .B(n483), .C(n267), .Y(o_dacv[90]) );
  OAI21BBX1 U367 ( .A(N1351), .B(n482), .C(n268), .Y(o_dacv[82]) );
  OAI21BBX1 U368 ( .A(N1395), .B(n486), .C(n281), .Y(o_dacv[114]) );
  OAI21BBX1 U369 ( .A(N1373), .B(n484), .C(n266), .Y(o_dacv[98]) );
  OAI21BBX1 U370 ( .A(N1384), .B(n485), .C(n282), .Y(o_dacv[106]) );
  OAI21BBX1 U371 ( .A(N1361), .B(n483), .C(n267), .Y(o_dacv[89]) );
  OAI21BBX1 U372 ( .A(N1350), .B(n482), .C(n268), .Y(o_dacv[81]) );
  OAI21BBX1 U373 ( .A(N1394), .B(n486), .C(n281), .Y(o_dacv[113]) );
  OAI21BBX1 U374 ( .A(N1372), .B(n484), .C(n266), .Y(o_dacv[97]) );
  OAI21BBX1 U375 ( .A(N1383), .B(n485), .C(n282), .Y(o_dacv[105]) );
  AO21X1 U376 ( .B(N1264), .C(n462), .A(n461), .Y(o_dacv[19]) );
  OAI21BBX1 U377 ( .A(N1386), .B(n485), .C(n282), .Y(o_dacv[108]) );
  AO21X1 U378 ( .B(N1262), .C(n462), .A(n461), .Y(o_dacv[17]) );
  AO21X1 U379 ( .B(N1263), .C(n462), .A(n461), .Y(o_dacv[18]) );
  AO21X1 U380 ( .B(N1268), .C(n462), .A(n461), .Y(o_dacv[23]) );
  INVX1 U381 ( .A(N1269), .Y(n462) );
  NOR21XL U382 ( .B(n223), .A(n243), .Y(n245) );
  GEN2XL U383 ( .D(n251), .E(n252), .C(n515), .B(n517), .A(n253), .Y(n246) );
  INVX1 U384 ( .A(n256), .Y(n515) );
  AOI21BBXL U385 ( .B(n249), .C(n250), .A(n517), .Y(n253) );
  GEN2XL U386 ( .D(n210), .E(n525), .C(n206), .B(n526), .A(n513), .Y(o_smpl[1]) );
  NAND3X1 U387 ( .A(n523), .B(n524), .C(n212), .Y(n210) );
  NAND21X1 U388 ( .B(n208), .A(n214), .Y(n211) );
  AND2X1 U389 ( .A(n254), .B(n252), .Y(n259) );
  OAI211X1 U390 ( .C(n246), .D(n518), .A(n247), .B(n517), .Y(n243) );
  INVX1 U391 ( .A(n140), .Y(n137) );
  AOI21X1 U392 ( .B(n223), .C(n227), .A(n514), .Y(n241) );
  OAI21BBX1 U393 ( .A(n251), .B(n254), .C(n255), .Y(n247) );
  OAI21BBX1 U394 ( .A(n231), .B(n226), .C(n232), .Y(n218) );
  OAI21X1 U395 ( .B(n239), .C(n229), .A(n240), .Y(n231) );
  OAI211X1 U396 ( .C(n216), .D(n524), .A(n218), .B(n523), .Y(n213) );
  OAI21X1 U397 ( .B(n241), .C(n229), .A(n233), .Y(n237) );
  NOR2X1 U398 ( .A(n525), .B(n214), .Y(n206) );
  NOR2X1 U399 ( .A(n213), .B(n204), .Y(n214) );
  INVX1 U400 ( .A(n258), .Y(n516) );
  NAND2X1 U401 ( .A(n245), .B(n519), .Y(n244) );
  NAND2X1 U402 ( .A(n230), .B(n247), .Y(n249) );
  NAND2X1 U403 ( .A(n238), .B(n521), .Y(n232) );
  INVX1 U404 ( .A(n236), .Y(n514) );
  INVX1 U405 ( .A(n209), .Y(n513) );
  INVX1 U406 ( .A(n140), .Y(n136) );
  INVX1 U407 ( .A(n139), .Y(n135) );
  INVX1 U408 ( .A(n139), .Y(r_adofs[7]) );
  NAND2X1 U409 ( .A(n233), .B(n234), .Y(n219) );
  GEN2XL U410 ( .D(n235), .E(n518), .C(n520), .B(n236), .A(n229), .Y(n234) );
  INVX1 U411 ( .A(n227), .Y(n520) );
  OAI21X1 U412 ( .B(n121), .C(n149), .A(n491), .Y(updlsb) );
  INVX1 U413 ( .A(n226), .Y(n522) );
  INVX1 U414 ( .A(n185), .Y(auto_sar) );
  NAND21X1 U415 ( .B(n101), .A(n89), .Y(n185) );
  INVX1 U416 ( .A(n159), .Y(n101) );
  NAND42X1 U417 ( .C(cs_ptr[3]), .D(n131), .A(tochg), .B(n528), .Y(n527) );
  INVX1 U418 ( .A(n149), .Y(n63) );
  NAND2X1 U419 ( .A(n128), .B(tochg), .Y(n528) );
  NAND2X1 U420 ( .A(n263), .B(n264), .Y(o_intr) );
  NOR4XL U421 ( .A(r_irq[7]), .B(r_irq[6]), .C(r_irq[5]), .D(r_irq[4]), .Y(
        n264) );
  NAND2X1 U422 ( .A(o_dactl[0]), .B(n89), .Y(n379) );
  NOR2X1 U423 ( .A(n150), .B(n494), .Y(updcmp) );
  XNOR2XL U424 ( .A(n89), .B(n94), .Y(n150) );
  AOI21X1 U425 ( .B(n159), .C(n160), .A(n494), .Y(sar_nxt) );
  NAND2X1 U426 ( .A(n94), .B(n89), .Y(n160) );
  NAND3X1 U427 ( .A(n525), .B(n526), .C(n204), .Y(o_smpl[4]) );
  AO21X1 U428 ( .B(N1251), .C(n459), .A(n458), .Y(o_dacv[9]) );
  AO21X1 U429 ( .B(N1250), .C(n459), .A(n458), .Y(o_dacv[8]) );
  AO21X1 U430 ( .B(N1254), .C(n459), .A(n458), .Y(o_dacv[12]) );
  AO21X1 U431 ( .B(N1257), .C(n459), .A(n458), .Y(o_dacv[15]) );
  AO21X1 U432 ( .B(N1311), .C(n474), .A(n473), .Y(o_dacv[54]) );
  AO21X1 U433 ( .B(N1310), .C(n474), .A(n473), .Y(o_dacv[53]) );
  AO21X1 U434 ( .B(N1278), .C(n465), .A(n464), .Y(o_dacv[30]) );
  AO21X1 U435 ( .B(N1277), .C(n465), .A(n464), .Y(o_dacv[29]) );
  AO21X1 U436 ( .B(N1279), .C(n465), .A(n464), .Y(o_dacv[31]) );
  AND2XL U437 ( .A(ps_ptr[4]), .B(r_sar_en[16]), .Y(n403) );
  AO21X1 U438 ( .B(N1312), .C(n474), .A(n473), .Y(o_dacv[55]) );
  AO21X1 U439 ( .B(N1305), .C(n474), .A(n473), .Y(o_dacv[48]) );
  AO21X1 U440 ( .B(N1308), .C(n474), .A(n473), .Y(o_dacv[51]) );
  AO21X1 U441 ( .B(N1307), .C(n474), .A(n473), .Y(o_dacv[50]) );
  AO21X1 U442 ( .B(N1317), .C(n477), .A(n476), .Y(o_dacv[57]) );
  AO21X1 U443 ( .B(N1319), .C(n477), .A(n476), .Y(o_dacv[59]) );
  AO21X1 U444 ( .B(N1316), .C(n477), .A(n476), .Y(o_dacv[56]) );
  AO21X1 U445 ( .B(N1318), .C(n477), .A(n476), .Y(o_dacv[58]) );
  AO21X1 U446 ( .B(N1323), .C(n477), .A(n476), .Y(o_dacv[63]) );
  AO2222X1 U447 ( .A(r_dac_en[9]), .B(n409), .C(r_dac_en[11]), .D(n408), .E(
        r_dac_en[13]), .F(n407), .G(r_dac_en[15]), .H(n406), .Y(n393) );
  AO21X1 U448 ( .B(N1261), .C(n462), .A(n461), .Y(o_dacv[16]) );
  AO21X1 U449 ( .B(N1283), .C(n468), .A(n467), .Y(o_dacv[32]) );
  AO21X1 U450 ( .B(N1272), .C(n465), .A(n464), .Y(o_dacv[24]) );
  AO21X1 U451 ( .B(N1255), .C(n459), .A(n458), .Y(o_dacv[13]) );
  AO21X1 U452 ( .B(N1252), .C(n459), .A(n458), .Y(o_dacv[10]) );
  AO21X1 U453 ( .B(N1256), .C(n459), .A(n458), .Y(o_dacv[14]) );
  AND2XL U454 ( .A(ps_ptr[4]), .B(r_dac_en[17]), .Y(n396) );
  NAND21X1 U455 ( .B(n198), .A(n197), .Y(n265) );
  NAND21X1 U456 ( .B(n433), .A(r_sar_en[15]), .Y(n194) );
  NOR43XL U457 ( .B(n190), .C(n189), .D(n188), .A(n187), .Y(n272) );
  NAND21X1 U458 ( .B(n445), .A(r_sar_en[5]), .Y(n190) );
  NAND21X1 U459 ( .B(n444), .A(r_sar_en[6]), .Y(n188) );
  NAND21X1 U460 ( .B(n447), .A(r_sar_en[4]), .Y(n189) );
  NAND21X1 U461 ( .B(n434), .A(r_sar_en[14]), .Y(n196) );
  NAND21X1 U462 ( .B(n435), .A(r_sar_en[13]), .Y(n195) );
  OAI21BBX1 U463 ( .A(N1422), .B(n488), .C(n279), .Y(o_dacv[135]) );
  OAI21BBX1 U464 ( .A(N1334), .B(n480), .C(n271), .Y(o_dacv[71]) );
  OAI21BBX1 U465 ( .A(N1345), .B(n481), .C(n270), .Y(o_dacv[79]) );
  OAI21BBX1 U466 ( .A(N1411), .B(n487), .C(n280), .Y(o_dacv[127]) );
  OAI21BBX1 U467 ( .A(N1433), .B(n489), .C(n278), .Y(o_dacv[143]) );
  AO21X1 U468 ( .B(N1239), .C(n456), .A(n455), .Y(o_dacv[0]) );
  AO21X1 U469 ( .B(N1294), .C(n471), .A(n470), .Y(o_dacv[40]) );
  NAND2X1 U470 ( .A(N1434), .B(n139), .Y(n278) );
  NAND2X1 U471 ( .A(N1346), .B(n139), .Y(n270) );
  NAND2X1 U472 ( .A(N1335), .B(n140), .Y(n271) );
  NAND2X1 U473 ( .A(N1368), .B(n140), .Y(n267) );
  NAND2X1 U474 ( .A(N1357), .B(n139), .Y(n268) );
  OAI21BBX1 U475 ( .A(N1420), .B(n488), .C(n279), .Y(o_dacv[133]) );
  OAI21BBX1 U476 ( .A(N1421), .B(n488), .C(n279), .Y(o_dacv[134]) );
  OAI21BBX1 U477 ( .A(N1415), .B(n488), .C(n279), .Y(o_dacv[128]) );
  OAI21BBX1 U478 ( .A(N1332), .B(n480), .C(n271), .Y(o_dacv[69]) );
  OAI21BBX1 U479 ( .A(N1409), .B(n487), .C(n280), .Y(o_dacv[125]) );
  OAI21BBX1 U480 ( .A(N1333), .B(n480), .C(n271), .Y(o_dacv[70]) );
  OAI21BBX1 U481 ( .A(N1410), .B(n487), .C(n280), .Y(o_dacv[126]) );
  OAI21BBX1 U482 ( .A(N1331), .B(n480), .C(n271), .Y(o_dacv[68]) );
  OAI21BBX1 U483 ( .A(N1408), .B(n487), .C(n280), .Y(o_dacv[124]) );
  OAI21BBX1 U484 ( .A(N1327), .B(n480), .C(n271), .Y(o_dacv[64]) );
  OAI21BBX1 U485 ( .A(N1404), .B(n487), .C(n280), .Y(o_dacv[120]) );
  OAI21BBX1 U486 ( .A(N1330), .B(n480), .C(n271), .Y(o_dacv[67]) );
  OAI21BBX1 U487 ( .A(N1407), .B(n487), .C(n280), .Y(o_dacv[123]) );
  OAI21BBX1 U488 ( .A(N1329), .B(n480), .C(n271), .Y(o_dacv[66]) );
  OAI21BBX1 U489 ( .A(N1328), .B(n480), .C(n271), .Y(o_dacv[65]) );
  OAI21BBX1 U490 ( .A(N1406), .B(n487), .C(n280), .Y(o_dacv[122]) );
  OAI21BBX1 U491 ( .A(N1405), .B(n487), .C(n280), .Y(o_dacv[121]) );
  OAI21BBX1 U492 ( .A(N1343), .B(n481), .C(n270), .Y(o_dacv[77]) );
  OAI21BBX1 U493 ( .A(N1344), .B(n481), .C(n270), .Y(o_dacv[78]) );
  OAI21BBX1 U494 ( .A(N1342), .B(n481), .C(n270), .Y(o_dacv[76]) );
  OAI21BBX1 U495 ( .A(N1338), .B(n481), .C(n270), .Y(o_dacv[72]) );
  OAI21BBX1 U496 ( .A(N1341), .B(n481), .C(n270), .Y(o_dacv[75]) );
  OAI21BBX1 U497 ( .A(N1340), .B(n481), .C(n270), .Y(o_dacv[74]) );
  OAI21BBX1 U498 ( .A(N1339), .B(n481), .C(n270), .Y(o_dacv[73]) );
  OAI21BBX1 U499 ( .A(N1431), .B(n489), .C(n278), .Y(o_dacv[141]) );
  OAI21BBX1 U500 ( .A(N1432), .B(n489), .C(n278), .Y(o_dacv[142]) );
  OAI21BBX1 U501 ( .A(N1426), .B(n489), .C(n278), .Y(o_dacv[136]) );
  MUX2AXL U502 ( .D0(r_rpt_v[6]), .D1(n24), .S(n121), .Y(n425) );
  OAI21BBX1 U503 ( .A(N1430), .B(n489), .C(n278), .Y(o_dacv[140]) );
  OAI21BBX1 U504 ( .A(N1419), .B(n488), .C(n279), .Y(o_dacv[132]) );
  OAI21BBX1 U505 ( .A(N1429), .B(n489), .C(n278), .Y(o_dacv[139]) );
  OAI21BBX1 U506 ( .A(N1418), .B(n488), .C(n279), .Y(o_dacv[131]) );
  OAI21BBX1 U507 ( .A(N1428), .B(n489), .C(n278), .Y(o_dacv[138]) );
  OAI21BBX1 U508 ( .A(N1427), .B(n489), .C(n278), .Y(o_dacv[137]) );
  OAI21BBX1 U509 ( .A(N1417), .B(n488), .C(n279), .Y(o_dacv[130]) );
  OAI21BBX1 U510 ( .A(N1416), .B(n488), .C(n279), .Y(o_dacv[129]) );
  OAI21BBX1 U511 ( .A(N1360), .B(n483), .C(n267), .Y(o_dacv[88]) );
  OAI21BBX1 U512 ( .A(N1349), .B(n482), .C(n268), .Y(o_dacv[80]) );
  OAI21BBX1 U513 ( .A(N1393), .B(n486), .C(n281), .Y(o_dacv[112]) );
  OAI21BBX1 U514 ( .A(N1371), .B(n484), .C(n266), .Y(o_dacv[96]) );
  ENOX1 U515 ( .A(n492), .B(n478), .C(r_rpt_v[9]), .D(n492), .Y(wda[7]) );
  ENOX1 U516 ( .A(n479), .B(n492), .C(r_rpt_v[8]), .D(n492), .Y(wda[6]) );
  MUX2AXL U517 ( .D0(r_rpt_v[2]), .D1(n429), .S(n121), .Y(n430) );
  MUX2AXL U518 ( .D0(r_rpt_v[5]), .D1(n426), .S(n121), .Y(n427) );
  MUX2AXL U519 ( .D0(r_rpt_v[4]), .D1(n20), .S(n121), .Y(n428) );
  MUX2AXL U520 ( .D0(r_rpt_v[7]), .D1(n27), .S(n121), .Y(n424) );
  INVX1 U521 ( .A(n460), .Y(n461) );
  NAND21X1 U522 ( .B(r_isofs[7]), .A(N1269), .Y(n460) );
  ENOX1 U523 ( .A(n479), .B(n491), .C(n491), .D(x_daclsb[5]), .Y(wdlsb[5]) );
  OAI21BBX1 U524 ( .A(N1382), .B(n485), .C(n282), .Y(o_dacv[104]) );
  XNOR2XL U525 ( .A(pos_dacis[1]), .B(pos_dacis[0]), .Y(n258) );
  AOI22AXL U526 ( .A(n255), .B(pos_dacis[5]), .D(n259), .C(pos_dacis[4]), .Y(
        n256) );
  AOI21BBXL U527 ( .B(n224), .C(n522), .A(n225), .Y(n212) );
  AOI211X1 U528 ( .C(n227), .D(n228), .A(n229), .B(n514), .Y(n224) );
  NAND32X1 U529 ( .B(n230), .C(pos_dacis[6]), .A(n518), .Y(n228) );
  GEN2XL U530 ( .D(n205), .E(n525), .C(n206), .B(n526), .A(n513), .Y(o_smpl[3]) );
  NAND42X1 U531 ( .C(pos_dacis[13]), .D(pos_dacis[14]), .A(n207), .B(n524), 
        .Y(n205) );
  AOI21BBXL U532 ( .B(pos_dacis[16]), .C(n215), .A(n206), .Y(n208) );
  NOR4XL U533 ( .A(pos_dacis[15]), .B(pos_dacis[14]), .C(n522), .D(n219), .Y(
        n215) );
  EORX1 U534 ( .A(n244), .B(pos_dacis[9]), .C(n245), .D(n519), .Y(n236) );
  NAND21X1 U535 ( .B(pos_dacis[4]), .A(n259), .Y(n255) );
  NAND21X1 U536 ( .B(pos_dacis[10]), .A(n242), .Y(n240) );
  ENOX1 U537 ( .A(n238), .B(n521), .C(n232), .D(pos_dacis[13]), .Y(n225) );
  OAI21X1 U538 ( .B(pos_dacis[3]), .C(n260), .A(n261), .Y(n252) );
  OAI21X1 U539 ( .B(n260), .C(n262), .A(pos_dacis[3]), .Y(n261) );
  EORX1 U540 ( .A(n262), .B(pos_dacis[2]), .C(pos_dacis[2]), .D(n516), .Y(n260) );
  NAND21X1 U541 ( .B(pos_dacis[0]), .A(n258), .Y(n262) );
  OAI22X1 U542 ( .A(pos_dacis[14]), .B(n220), .C(n221), .D(n523), .Y(n216) );
  AOI21X1 U543 ( .B(n226), .C(n237), .A(n225), .Y(n220) );
  NOR42XL U544 ( .C(n219), .D(n218), .A(n212), .B(n207), .Y(n221) );
  AOI22AXL U545 ( .A(n240), .B(pos_dacis[11]), .D(n242), .C(pos_dacis[10]), 
        .Y(n233) );
  EORX1 U546 ( .A(n524), .B(n216), .C(n217), .D(n524), .Y(n204) );
  NOR32XL U547 ( .B(n216), .C(n218), .A(pos_dacis[14]), .Y(n217) );
  NAND2X1 U548 ( .A(pos_dacis[17]), .B(n211), .Y(n209) );
  OAI21BBX1 U549 ( .A(n518), .B(n246), .C(n248), .Y(n223) );
  OAI31XL U550 ( .A(n249), .B(pos_dacis[6]), .C(n235), .D(pos_dacis[7]), .Y(
        n248) );
  OAI31XL U551 ( .A(n213), .B(pos_dacis[17]), .C(pos_dacis[16]), .D(n211), .Y(
        o_smpl[0]) );
  OAI21X1 U552 ( .B(pos_dacis[17]), .C(n208), .A(n209), .Y(o_smpl[2]) );
  INVX1 U553 ( .A(n534), .Y(n140) );
  NAND2X1 U554 ( .A(n256), .B(n257), .Y(n230) );
  OAI31XL U555 ( .A(n258), .B(pos_dacis[3]), .C(pos_dacis[2]), .D(n251), .Y(
        n257) );
  NOR32XL U556 ( .B(n250), .C(n517), .A(pos_dacis[5]), .Y(n235) );
  AOI211X1 U557 ( .C(n516), .D(pos_dacis[3]), .A(pos_dacis[0]), .B(
        pos_dacis[2]), .Y(n254) );
  INVX1 U558 ( .A(n534), .Y(n139) );
  NOR2X1 U559 ( .A(n252), .B(pos_dacis[4]), .Y(n250) );
  NOR32XL U560 ( .B(n193), .C(n192), .A(n191), .Y(n269) );
  NAND2X1 U561 ( .A(r_sar_en[3]), .B(dacv_wr[3]), .Y(n192) );
  NAND2X1 U562 ( .A(r_sar_en[2]), .B(dacv_wr[2]), .Y(n193) );
  AO22X1 U563 ( .A(r_sar_en[0]), .B(dacv_wr[0]), .C(r_sar_en[1]), .D(
        dacv_wr[1]), .Y(n191) );
  NOR42XL U564 ( .C(n519), .D(n222), .A(pos_dacis[12]), .B(pos_dacis[9]), .Y(
        n207) );
  NOR3XL U565 ( .A(n223), .B(pos_dacis[11]), .C(pos_dacis[10]), .Y(n222) );
  NOR2X1 U566 ( .A(pos_dacis[4]), .B(pos_dacis[5]), .Y(n251) );
  INVX1 U567 ( .A(pos_dacis[6]), .Y(n517) );
  NOR21XL U568 ( .B(app_dacis[11]), .A(r_comp_opt[0]), .Y(o_daci_sel[11]) );
  NOR21XL U569 ( .B(app_dacis[6]), .A(n69), .Y(o_daci_sel[6]) );
  NOR21XL U570 ( .B(app_dacis[7]), .A(n69), .Y(o_daci_sel[7]) );
  NOR21XL U571 ( .B(app_dacis[16]), .A(n69), .Y(o_daci_sel[16]) );
  NOR21XL U572 ( .B(app_dacis[0]), .A(n69), .Y(o_daci_sel[0]) );
  INVX1 U573 ( .A(pos_dacis[7]), .Y(n518) );
  NOR21XL U574 ( .B(app_dacis[14]), .A(n69), .Y(o_daci_sel[14]) );
  NOR21XL U575 ( .B(app_dacis[12]), .A(r_comp_opt[0]), .Y(o_daci_sel[12]) );
  NOR21XL U576 ( .B(app_dacis[15]), .A(n69), .Y(o_daci_sel[15]) );
  NOR21XL U577 ( .B(app_dacis[5]), .A(n69), .Y(o_daci_sel[5]) );
  NOR21XL U578 ( .B(app_dacis[17]), .A(n69), .Y(o_daci_sel[17]) );
  NOR21XL U579 ( .B(app_dacis[2]), .A(r_comp_opt[0]), .Y(o_daci_sel[2]) );
  NOR21XL U580 ( .B(app_dacis[3]), .A(r_comp_opt[0]), .Y(o_daci_sel[3]) );
  NOR21XL U581 ( .B(app_dacis[13]), .A(r_comp_opt[0]), .Y(o_daci_sel[13]) );
  NOR21XL U582 ( .B(app_dacis[10]), .A(r_comp_opt[0]), .Y(o_daci_sel[10]) );
  NOR21XL U583 ( .B(app_dacis[8]), .A(r_comp_opt[0]), .Y(o_daci_sel[8]) );
  NOR21XL U584 ( .B(app_dacis[4]), .A(n69), .Y(o_daci_sel[4]) );
  NOR21XL U585 ( .B(app_dacis[1]), .A(n69), .Y(o_daci_sel[1]) );
  NOR21XL U586 ( .B(app_dacis[9]), .A(r_comp_opt[0]), .Y(o_daci_sel[9]) );
  NOR2X1 U587 ( .A(pos_dacis[8]), .B(pos_dacis[9]), .Y(n227) );
  INVX1 U588 ( .A(pos_dacis[8]), .Y(n519) );
  OR2X1 U589 ( .A(pos_dacis[11]), .B(pos_dacis[10]), .Y(n229) );
  NOR2X1 U590 ( .A(pos_dacis[12]), .B(pos_dacis[13]), .Y(n226) );
  INVX1 U591 ( .A(pos_dacis[12]), .Y(n521) );
  INVX1 U592 ( .A(pos_dacis[14]), .Y(n523) );
  INVX1 U593 ( .A(pos_dacis[15]), .Y(n524) );
  INVX1 U594 ( .A(pos_dacis[16]), .Y(n525) );
  INVX1 U595 ( .A(pos_dacis[17]), .Y(n526) );
  NAND42X1 U596 ( .C(r_dac_en[4]), .D(n184), .A(n183), .B(n182), .Y(n159) );
  NOR43XL U597 ( .B(n181), .C(n180), .D(n179), .A(n178), .Y(n182) );
  NAND21X1 U598 ( .B(r_dac_en[2]), .A(n176), .Y(n184) );
  NOR32XL U599 ( .B(n93), .C(n92), .A(n177), .Y(n183) );
  MUX4X1 U600 ( .D0(r_sar_en[2]), .D1(r_sar_en[3]), .D2(r_sar_en[10]), .D3(
        r_sar_en[11]), .S0(n117), .S1(n115), .Y(n105) );
  MUX4X1 U601 ( .D0(r_sar_en[4]), .D1(r_sar_en[5]), .D2(r_sar_en[12]), .D3(
        r_sar_en[13]), .S0(n117), .S1(n115), .Y(n106) );
  MUX4X1 U602 ( .D0(r_sar_en[0]), .D1(r_sar_en[1]), .D2(r_sar_en[8]), .D3(
        r_sar_en[9]), .S0(n117), .S1(n115), .Y(n107) );
  MUX4X1 U603 ( .D0(r_sar_en[6]), .D1(r_sar_en[7]), .D2(r_sar_en[14]), .D3(
        r_sar_en[15]), .S0(n117), .S1(n115), .Y(n104) );
  INVX1 U604 ( .A(r_dac_en[3]), .Y(n176) );
  OR4X1 U605 ( .A(r_dac_en[5]), .B(r_dac_en[6]), .C(r_dac_en[11]), .D(
        r_dac_en[10]), .Y(n178) );
  INVX1 U606 ( .A(r_dac_en[14]), .Y(n179) );
  INVX1 U607 ( .A(r_dac_en[13]), .Y(n181) );
  INVX1 U608 ( .A(r_dac_en[12]), .Y(n180) );
  MUX2BXL U609 ( .D0(n90), .D1(n91), .S(n131), .Y(n89) );
  MUX4X1 U610 ( .D0(n107), .D1(n105), .D2(n106), .D3(n104), .S0(n126), .S1(
        n128), .Y(n90) );
  MUX2IX1 U611 ( .D0(r_sar_en[16]), .D1(r_sar_en[17]), .S(n116), .Y(n91) );
  OR2X1 U612 ( .A(r_dac_en[0]), .B(r_dac_en[1]), .Y(n177) );
  NOR3XL U613 ( .A(r_dac_en[15]), .B(r_dac_en[16]), .C(r_dac_en[17]), .Y(n92)
         );
  NOR3XL U614 ( .A(r_dac_en[7]), .B(r_dac_en[8]), .C(r_dac_en[9]), .Y(n93) );
  MUX4X1 U615 ( .D0(n112), .D1(n110), .D2(n111), .D3(n109), .S0(n126), .S1(
        n128), .Y(n113) );
  MUX4X1 U616 ( .D0(o_dat[4]), .D1(o_dat[5]), .D2(o_dat[12]), .D3(o_dat[13]), 
        .S0(n116), .S1(n115), .Y(n111) );
  MUX4X1 U617 ( .D0(o_dat[6]), .D1(o_dat[7]), .D2(o_dat[14]), .D3(o_dat[15]), 
        .S0(n117), .S1(n115), .Y(n109) );
  MUX4X1 U618 ( .D0(o_dat[2]), .D1(o_dat[3]), .D2(o_dat[10]), .D3(o_dat[11]), 
        .S0(n116), .S1(n115), .Y(n110) );
  MUX4X1 U619 ( .D0(o_dat[0]), .D1(o_dat[1]), .D2(o_dat[8]), .D3(o_dat[9]), 
        .S0(n117), .S1(n115), .Y(n112) );
  NOR42XL U620 ( .C(o_dactl[1]), .D(dacyc_done), .A(n89), .B(n152), .Y(tochg)
         );
  XNOR2XL U621 ( .A(syn_comp[1]), .B(N859), .Y(n152) );
  MUX2X1 U622 ( .D0(n113), .D1(n108), .S(n131), .Y(N859) );
  MUX2X1 U623 ( .D0(o_dat[16]), .D1(o_dat[17]), .S(n116), .Y(n108) );
  XNOR2XL U624 ( .A(n127), .B(x_daclsb[4]), .Y(n203) );
  NAND4X1 U625 ( .A(o_dactl[6]), .B(n199), .C(n200), .D(n201), .Y(n149) );
  NOR2X1 U626 ( .A(n202), .B(n203), .Y(n201) );
  XNOR2XL U627 ( .A(x_daclsb[3]), .B(n124), .Y(n200) );
  XNOR2XL U628 ( .A(n129), .B(x_daclsb[5]), .Y(n202) );
  NOR4XL U629 ( .A(r_irq[3]), .B(r_irq[2]), .C(r_irq[1]), .D(r_irq[0]), .Y(
        n263) );
  AO222X1 U630 ( .A(n283), .B(n364), .C(n285), .D(n365), .E(r_dac1v[2]), .F(
        n493), .Y(o_dac1[2]) );
  NAND4X1 U631 ( .A(n370), .B(n371), .C(n372), .D(n373), .Y(n364) );
  NAND4X1 U632 ( .A(n366), .B(n367), .C(n368), .D(n369), .Y(n365) );
  AOI22X1 U633 ( .A(r_dacvs[8]), .B(n43), .C(r_dacvs[136]), .D(n68), .Y(n370)
         );
  AO222X1 U634 ( .A(n283), .B(n354), .C(n285), .D(n355), .E(r_dac1v[3]), .F(
        n493), .Y(o_dac1[3]) );
  NAND4X1 U635 ( .A(n360), .B(n361), .C(n362), .D(n363), .Y(n354) );
  NAND4X1 U636 ( .A(n356), .B(n357), .C(n358), .D(n359), .Y(n355) );
  AOI22X1 U637 ( .A(r_dacvs[9]), .B(n43), .C(r_dacvs[137]), .D(n68), .Y(n360)
         );
  AO222X1 U638 ( .A(n283), .B(n344), .C(n285), .D(n345), .E(r_dac1v[4]), .F(
        n493), .Y(o_dac1[4]) );
  NAND4X1 U639 ( .A(n350), .B(n351), .C(n352), .D(n353), .Y(n344) );
  NAND4X1 U640 ( .A(n346), .B(n347), .C(n348), .D(n349), .Y(n345) );
  AOI22X1 U641 ( .A(r_dacvs[10]), .B(n43), .C(r_dacvs[138]), .D(n68), .Y(n350)
         );
  AO222X1 U642 ( .A(n283), .B(n324), .C(n285), .D(n325), .E(r_dac1v[6]), .F(
        n493), .Y(o_dac1[6]) );
  NAND4X1 U643 ( .A(n330), .B(n331), .C(n332), .D(n333), .Y(n324) );
  NAND4X1 U644 ( .A(n326), .B(n327), .C(n328), .D(n329), .Y(n325) );
  AOI22X1 U645 ( .A(r_dacvs[12]), .B(n42), .C(r_dacvs[140]), .D(n299), .Y(n330) );
  AO222X1 U646 ( .A(n283), .B(n314), .C(n285), .D(n315), .E(r_dac1v[7]), .F(
        n493), .Y(o_dac1[7]) );
  NAND4X1 U647 ( .A(n320), .B(n321), .C(n322), .D(n323), .Y(n314) );
  NAND4X1 U648 ( .A(n316), .B(n317), .C(n318), .D(n319), .Y(n315) );
  AOI22X1 U649 ( .A(r_dacvs[13]), .B(n43), .C(r_dacvs[141]), .D(n68), .Y(n320)
         );
  AO222X1 U650 ( .A(n283), .B(n304), .C(n285), .D(n305), .E(r_dac1v[8]), .F(
        n493), .Y(o_dac1[8]) );
  NAND4X1 U651 ( .A(n310), .B(n311), .C(n312), .D(n313), .Y(n304) );
  NAND4X1 U652 ( .A(n306), .B(n307), .C(n308), .D(n309), .Y(n305) );
  AOI22X1 U653 ( .A(r_dacvs[14]), .B(n43), .C(r_dacvs[142]), .D(n299), .Y(n310) );
  AO222X1 U654 ( .A(n283), .B(n284), .C(n285), .D(n286), .E(r_dac1v[9]), .F(
        n493), .Y(o_dac1[9]) );
  NAND4X1 U655 ( .A(n300), .B(n301), .C(n302), .D(n303), .Y(n284) );
  NAND4X1 U656 ( .A(n287), .B(n288), .C(n289), .D(n290), .Y(n286) );
  AOI22X1 U657 ( .A(r_dacvs[15]), .B(n42), .C(r_dacvs[143]), .D(n299), .Y(n300) );
  AO222X1 U658 ( .A(n283), .B(n334), .C(n285), .D(n335), .E(r_dac1v[5]), .F(
        n493), .Y(o_dac1[5]) );
  NAND4X1 U659 ( .A(n340), .B(n341), .C(n342), .D(n343), .Y(n334) );
  NAND4X1 U660 ( .A(n336), .B(n337), .C(n338), .D(n339), .Y(n335) );
  AOI22X1 U661 ( .A(r_dacvs[11]), .B(n43), .C(r_dacvs[139]), .D(n299), .Y(n340) );
  AO22X1 U662 ( .A(r_dac1v[0]), .B(n493), .C(x_daclsb[0]), .D(n379), .Y(
        o_dac1[0]) );
  AO22X1 U663 ( .A(r_dac1v[1]), .B(n493), .C(x_daclsb[1]), .D(n379), .Y(
        o_dac1[1]) );
  MUX4X1 U664 ( .D0(r_dac_en[2]), .D1(r_dac_en[3]), .D2(r_dac_en[10]), .D3(
        r_dac_en[11]), .S0(n117), .S1(n114), .Y(n100) );
  MUX4X1 U665 ( .D0(r_dac_en[0]), .D1(r_dac_en[1]), .D2(r_dac_en[8]), .D3(
        r_dac_en[9]), .S0(n117), .S1(n115), .Y(n103) );
  MUX4X1 U666 ( .D0(r_dac_en[4]), .D1(r_dac_en[5]), .D2(r_dac_en[12]), .D3(
        r_dac_en[13]), .S0(n117), .S1(n115), .Y(n102) );
  MUX4X1 U667 ( .D0(r_dac_en[6]), .D1(r_dac_en[7]), .D2(r_dac_en[14]), .D3(
        r_dac_en[15]), .S0(n117), .S1(n114), .Y(n97) );
  AOI222XL U668 ( .A(r_dacvs[115]), .B(n52), .C(r_dacvs[83]), .D(n59), .E(
        r_dacvs[99]), .F(n66), .Y(n339) );
  AOI222XL U669 ( .A(r_dacvs[123]), .B(n53), .C(r_dacvs[91]), .D(n60), .E(
        r_dacvs[107]), .F(n67), .Y(n343) );
  AOI222XL U670 ( .A(r_dacvs[116]), .B(n52), .C(r_dacvs[84]), .D(n59), .E(
        r_dacvs[100]), .F(n66), .Y(n329) );
  AOI222XL U671 ( .A(r_dacvs[124]), .B(n52), .C(r_dacvs[92]), .D(n59), .E(
        r_dacvs[108]), .F(n66), .Y(n333) );
  AOI222XL U672 ( .A(r_dacvs[118]), .B(n52), .C(r_dacvs[86]), .D(n59), .E(
        r_dacvs[102]), .F(n66), .Y(n309) );
  AOI222XL U673 ( .A(r_dacvs[126]), .B(n53), .C(r_dacvs[94]), .D(n60), .E(
        r_dacvs[110]), .F(n67), .Y(n313) );
  AOI222XL U674 ( .A(r_dacvs[119]), .B(n52), .C(r_dacvs[87]), .D(n59), .E(
        r_dacvs[103]), .F(n66), .Y(n290) );
  AOI222XL U675 ( .A(r_dacvs[127]), .B(n52), .C(r_dacvs[95]), .D(n59), .E(
        r_dacvs[111]), .F(n66), .Y(n303) );
  AOI22X1 U676 ( .A(r_dacvs[67]), .B(n46), .C(r_dacvs[19]), .D(n64), .Y(n338)
         );
  AOI22X1 U677 ( .A(r_dacvs[75]), .B(n47), .C(r_dacvs[27]), .D(n65), .Y(n342)
         );
  AOI22X1 U678 ( .A(r_dacvs[68]), .B(n46), .C(r_dacvs[20]), .D(n64), .Y(n328)
         );
  AOI22X1 U679 ( .A(r_dacvs[70]), .B(n46), .C(r_dacvs[22]), .D(n64), .Y(n308)
         );
  AOI22X1 U680 ( .A(r_dacvs[71]), .B(n46), .C(r_dacvs[23]), .D(n64), .Y(n289)
         );
  AOI22X1 U681 ( .A(r_dacvs[79]), .B(n46), .C(r_dacvs[31]), .D(n64), .Y(n302)
         );
  MUX2BXL U682 ( .D0(n95), .D1(n96), .S(n131), .Y(n94) );
  MUX4X1 U683 ( .D0(n103), .D1(n100), .D2(n102), .D3(n97), .S0(n126), .S1(n128), .Y(n95) );
  MUX2IX1 U684 ( .D0(r_dac_en[16]), .D1(r_dac_en[17]), .S(n116), .Y(n96) );
  AOI22X1 U685 ( .A(r_dacvs[35]), .B(n50), .C(r_dacvs[51]), .D(n57), .Y(n337)
         );
  AOI22X1 U686 ( .A(r_dacvs[36]), .B(n50), .C(r_dacvs[52]), .D(n57), .Y(n327)
         );
  AOI22X1 U687 ( .A(r_dacvs[38]), .B(n50), .C(r_dacvs[54]), .D(n57), .Y(n307)
         );
  AOI22X1 U688 ( .A(r_dacvs[39]), .B(n50), .C(r_dacvs[55]), .D(n57), .Y(n288)
         );
  AOI22X1 U689 ( .A(r_dacvs[3]), .B(n42), .C(r_dacvs[131]), .D(n299), .Y(n336)
         );
  AOI22X1 U690 ( .A(r_dacvs[4]), .B(n42), .C(r_dacvs[132]), .D(n299), .Y(n326)
         );
  AOI22X1 U691 ( .A(r_dacvs[7]), .B(n42), .C(r_dacvs[135]), .D(n299), .Y(n287)
         );
  AOI222XL U692 ( .A(r_dacvs[112]), .B(n53), .C(r_dacvs[80]), .D(n60), .E(
        r_dacvs[96]), .F(n67), .Y(n369) );
  AOI222XL U693 ( .A(r_dacvs[120]), .B(n53), .C(r_dacvs[88]), .D(n60), .E(
        r_dacvs[104]), .F(n67), .Y(n373) );
  AOI222XL U694 ( .A(r_dacvs[113]), .B(n53), .C(r_dacvs[81]), .D(n60), .E(
        r_dacvs[97]), .F(n67), .Y(n359) );
  AOI222XL U695 ( .A(r_dacvs[121]), .B(n53), .C(r_dacvs[89]), .D(n60), .E(
        r_dacvs[105]), .F(n67), .Y(n363) );
  AOI222XL U696 ( .A(r_dacvs[114]), .B(n53), .C(r_dacvs[82]), .D(n60), .E(
        r_dacvs[98]), .F(n67), .Y(n349) );
  AOI222XL U697 ( .A(r_dacvs[122]), .B(n53), .C(r_dacvs[90]), .D(n60), .E(
        r_dacvs[106]), .F(n67), .Y(n353) );
  AOI222XL U698 ( .A(r_dacvs[117]), .B(n53), .C(r_dacvs[85]), .D(n60), .E(
        r_dacvs[101]), .F(n67), .Y(n319) );
  AOI222XL U699 ( .A(r_dacvs[125]), .B(n53), .C(r_dacvs[93]), .D(n60), .E(
        r_dacvs[109]), .F(n67), .Y(n323) );
  AOI22X1 U700 ( .A(r_dacvs[64]), .B(n47), .C(r_dacvs[16]), .D(n65), .Y(n368)
         );
  AOI22X1 U701 ( .A(r_dacvs[72]), .B(n47), .C(r_dacvs[24]), .D(n65), .Y(n372)
         );
  AOI22X1 U702 ( .A(r_dacvs[65]), .B(n47), .C(r_dacvs[17]), .D(n65), .Y(n358)
         );
  AOI22X1 U703 ( .A(r_dacvs[73]), .B(n47), .C(r_dacvs[25]), .D(n65), .Y(n362)
         );
  AOI22X1 U704 ( .A(r_dacvs[66]), .B(n47), .C(r_dacvs[18]), .D(n65), .Y(n348)
         );
  AOI22X1 U705 ( .A(r_dacvs[74]), .B(n47), .C(r_dacvs[26]), .D(n65), .Y(n352)
         );
  AOI22X1 U706 ( .A(r_dacvs[76]), .B(n46), .C(r_dacvs[28]), .D(n64), .Y(n332)
         );
  AOI22X1 U707 ( .A(r_dacvs[69]), .B(n47), .C(r_dacvs[21]), .D(n65), .Y(n318)
         );
  AOI22X1 U708 ( .A(r_dacvs[77]), .B(n47), .C(r_dacvs[29]), .D(n65), .Y(n322)
         );
  AOI22X1 U709 ( .A(r_dacvs[78]), .B(n47), .C(r_dacvs[30]), .D(n65), .Y(n312)
         );
  AOI22X1 U710 ( .A(r_dacvs[32]), .B(n51), .C(r_dacvs[48]), .D(n58), .Y(n367)
         );
  AOI22X1 U711 ( .A(r_dacvs[40]), .B(n51), .C(r_dacvs[56]), .D(n58), .Y(n371)
         );
  AOI22X1 U712 ( .A(r_dacvs[33]), .B(n51), .C(r_dacvs[49]), .D(n58), .Y(n357)
         );
  AOI22X1 U713 ( .A(r_dacvs[41]), .B(n51), .C(r_dacvs[57]), .D(n58), .Y(n361)
         );
  AOI22X1 U714 ( .A(r_dacvs[34]), .B(n51), .C(r_dacvs[50]), .D(n58), .Y(n347)
         );
  AOI22X1 U715 ( .A(r_dacvs[42]), .B(n51), .C(r_dacvs[58]), .D(n58), .Y(n351)
         );
  AOI22X1 U716 ( .A(r_dacvs[43]), .B(n51), .C(r_dacvs[59]), .D(n58), .Y(n341)
         );
  AOI22X1 U717 ( .A(r_dacvs[44]), .B(n50), .C(r_dacvs[60]), .D(n57), .Y(n331)
         );
  AOI22X1 U718 ( .A(r_dacvs[37]), .B(n51), .C(r_dacvs[53]), .D(n58), .Y(n317)
         );
  AOI22X1 U719 ( .A(r_dacvs[45]), .B(n51), .C(r_dacvs[61]), .D(n58), .Y(n321)
         );
  AOI22X1 U720 ( .A(r_dacvs[46]), .B(n51), .C(r_dacvs[62]), .D(n58), .Y(n311)
         );
  AOI22X1 U721 ( .A(r_dacvs[47]), .B(n50), .C(r_dacvs[63]), .D(n57), .Y(n301)
         );
  AOI22X1 U722 ( .A(r_dacvs[0]), .B(n43), .C(r_dacvs[128]), .D(n299), .Y(n366)
         );
  AOI22X1 U723 ( .A(r_dacvs[1]), .B(n43), .C(r_dacvs[129]), .D(n68), .Y(n356)
         );
  AOI22X1 U724 ( .A(r_dacvs[2]), .B(n43), .C(r_dacvs[130]), .D(n68), .Y(n346)
         );
  AOI22X1 U725 ( .A(r_dacvs[5]), .B(n43), .C(r_dacvs[133]), .D(n68), .Y(n316)
         );
  AOI22X1 U726 ( .A(r_dacvs[6]), .B(n42), .C(r_dacvs[134]), .D(n299), .Y(n306)
         );
  INVX1 U727 ( .A(r_sar_en[17]), .Y(n404) );
  ENOX1 U728 ( .A(n502), .B(n134), .C(o_dat[2]), .D(n502), .Y(datcmp[2]) );
  ENOX1 U729 ( .A(n506), .B(n134), .C(o_dat[3]), .D(n506), .Y(datcmp[3]) );
  ENOX1 U730 ( .A(n498), .B(n134), .C(o_dat[4]), .D(n498), .Y(datcmp[4]) );
  ENOX1 U731 ( .A(n511), .B(n134), .C(o_dat[5]), .D(n511), .Y(datcmp[5]) );
  ENOX1 U732 ( .A(n503), .B(n134), .C(o_dat[6]), .D(n503), .Y(datcmp[6]) );
  ENOX1 U733 ( .A(n507), .B(n134), .C(o_dat[7]), .D(n507), .Y(datcmp[7]) );
  ENOX1 U734 ( .A(n499), .B(n134), .C(o_dat[8]), .D(n499), .Y(datcmp[8]) );
  ENOX1 U735 ( .A(n512), .B(n134), .C(o_dat[9]), .D(n512), .Y(datcmp[9]) );
  ENOX1 U736 ( .A(n495), .B(n133), .C(o_dat[0]), .D(n495), .Y(datcmp[0]) );
  ENOX1 U737 ( .A(n510), .B(n133), .C(o_dat[1]), .D(n510), .Y(datcmp[1]) );
  ENOX1 U738 ( .A(n500), .B(n133), .C(o_dat[10]), .D(n500), .Y(datcmp[10]) );
  ENOX1 U739 ( .A(n504), .B(n133), .C(o_dat[11]), .D(n504), .Y(datcmp[11]) );
  ENOX1 U740 ( .A(n496), .B(n133), .C(o_dat[12]), .D(n496), .Y(datcmp[12]) );
  ENOX1 U741 ( .A(n508), .B(n133), .C(o_dat[13]), .D(n508), .Y(datcmp[13]) );
  ENOX1 U742 ( .A(n501), .B(n133), .C(o_dat[14]), .D(n501), .Y(datcmp[14]) );
  ENOX1 U743 ( .A(n505), .B(n133), .C(o_dat[15]), .D(n505), .Y(datcmp[15]) );
  ENOX1 U744 ( .A(n497), .B(n133), .C(o_dat[16]), .D(n497), .Y(datcmp[16]) );
  ENOX1 U745 ( .A(n509), .B(n133), .C(o_dat[17]), .D(n509), .Y(datcmp[17]) );
  INVX1 U746 ( .A(syn_comp[1]), .Y(n133) );
  INVX1 U747 ( .A(syn_comp[1]), .Y(n134) );
  INVXL U748 ( .A(dacv_wr[10]), .Y(n439) );
  BUFXL U749 ( .A(r_wdat[0]), .Y(n118) );
  BUFXL U750 ( .A(r_wdat[0]), .Y(n119) );
  NAND21X2 U751 ( .B(n413), .A(n412), .Y(n414) );
  MUX2IX2 U752 ( .D0(n411), .D1(n410), .S(ps_ptr[3]), .Y(n412) );
  NAND21X2 U753 ( .B(n403), .A(n402), .Y(n415) );
  MUX2IX2 U754 ( .D0(n401), .D1(n400), .S(ps_ptr[3]), .Y(n402) );
  AO2222X1 U755 ( .A(n408), .B(r_sar_en[3]), .C(n405), .D(r_sar_en[1]), .E(
        n407), .F(r_sar_en[5]), .G(n406), .H(r_sar_en[7]), .Y(n411) );
  INVXL U756 ( .A(ps_ptr[4]), .Y(n382) );
  MUX2IX2 U757 ( .D0(n394), .D1(n393), .S(ps_ptr[3]), .Y(n395) );
  NAND21X2 U758 ( .B(n392), .A(n391), .Y(n398) );
  INVXL U759 ( .A(n98), .Y(n380) );
  NAND32X2 U760 ( .B(n101), .C(n19), .A(n98), .Y(n399) );
  INVXL U761 ( .A(n118), .Y(n429) );
  AND2XL U762 ( .A(n119), .B(r_wr[4]), .Y(clrsta[0]) );
  NAND6XL U763 ( .A(r_wdat[6]), .B(n119), .C(n277), .D(n20), .E(n426), .F(n27), 
        .Y(n276) );
  MUX2XL U764 ( .D0(n29), .D1(o_dactl[5]), .S(n380), .Y(ps_md4ch) );
  MUX2XL U765 ( .D0(n25), .D1(x_daclsb[3]), .S(n491), .Y(wdlsb[3]) );
  MUX2XL U766 ( .D0(n26), .D1(o_dactl[4]), .S(n380), .Y(ps_sample) );
  NOR32XL U767 ( .B(n101), .C(r_wdat[7]), .A(o_dactl[0]), .Y(n274) );
  NOR21XL U768 ( .B(n22), .A(n25), .Y(n275) );
  MUX2X1 U769 ( .D0(n28), .D1(x_daclsb[4]), .S(n491), .Y(wdlsb[4]) );
  NAND6XL U770 ( .A(n29), .B(r_wdat[3]), .C(n21), .D(n277), .E(n429), .F(n479), 
        .Y(n381) );
  MUX2X1 U771 ( .D0(n21), .D1(x_daclsb[2]), .S(n491), .Y(wdlsb[2]) );
  MUX2XL U772 ( .D0(n23), .D1(r_rpt_v[1]), .S(n491), .Y(wdlsb[1]) );
  MUX2XL U773 ( .D0(n118), .D1(r_rpt_v[0]), .S(n491), .Y(wdlsb[0]) );
  AO22XL U774 ( .A(dacv_wr[8]), .B(r_sar_en[8]), .C(dacv_wr[7]), .D(
        r_sar_en[7]), .Y(n187) );
  AO2222X1 U775 ( .A(n409), .B(r_sar_en[8]), .C(n408), .D(r_sar_en[10]), .E(
        n407), .F(r_sar_en[12]), .G(n406), .H(r_sar_en[14]), .Y(n400) );
  INVXL U776 ( .A(dacv_wr[14]), .Y(n434) );
  AO2222XL U777 ( .A(dacv_wr[10]), .B(r_sar_en[10]), .C(dacv_wr[11]), .D(
        r_sar_en[11]), .E(dacv_wr[9]), .F(r_sar_en[9]), .G(dacv_wr[12]), .H(
        r_sar_en[12]), .Y(n198) );
  INVXL U778 ( .A(dacv_wr[12]), .Y(n436) );
  AO2222X1 U779 ( .A(r_dac_en[2]), .B(n408), .C(r_dac_en[0]), .D(n405), .E(
        r_dac_en[4]), .F(n407), .G(r_dac_en[6]), .H(n406), .Y(n390) );
  INVX3 U780 ( .A(n385), .Y(n405) );
  NAND21X2 U781 ( .B(n396), .A(n395), .Y(n397) );
  MUX2IX2 U782 ( .D0(n398), .D1(n397), .S(ps_ptr[0]), .Y(n419) );
  AO2222X1 U783 ( .A(n408), .B(r_sar_en[2]), .C(n405), .D(r_sar_en[0]), .E(
        n407), .F(r_sar_en[4]), .G(n406), .H(r_sar_en[6]), .Y(n401) );
  NOR21XL U784 ( .B(ps_ptr[4]), .A(n404), .Y(n413) );
  AO2222X1 U785 ( .A(r_dac_en[3]), .B(n408), .C(r_dac_en[1]), .D(n405), .E(
        r_dac_en[5]), .F(n407), .G(r_dac_en[7]), .H(n406), .Y(n394) );
  NAND21XL U786 ( .B(n87), .A(n399), .Y(n417) );
  AO21X4 U787 ( .B(r_wr[0]), .C(n186), .A(n19), .Y(n98) );
  NAND21X4 U788 ( .B(ps_ptr[2]), .A(ps_ptr[1]), .Y(n383) );
  INVX8 U789 ( .A(n383), .Y(n408) );
endmodule


module dacmux_a0_DW01_add_17 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;

  wire   [8:1] carry;

  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  XOR2X1 U1 ( .A(B[8]), .B(carry[8]), .Y(SUM[8]) );
  AND2X1 U2 ( .A(A[0]), .B(B[0]), .Y(carry[1]) );
  XOR2XL U3 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
endmodule


module dacmux_a0_DW01_add_16 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;

  wire   [8:1] carry;

  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  XOR2X1 U1 ( .A(B[8]), .B(carry[8]), .Y(SUM[8]) );
  XOR2X1 U2 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
  AND2X1 U3 ( .A(A[0]), .B(B[0]), .Y(carry[1]) );
endmodule


module dacmux_a0_DW01_add_15 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;

  wire   [8:1] carry;

  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  XOR2X1 U1 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
  AND2X1 U2 ( .A(A[0]), .B(B[0]), .Y(carry[1]) );
  XOR2X1 U3 ( .A(B[8]), .B(carry[8]), .Y(SUM[8]) );
endmodule


module dacmux_a0_DW01_add_14 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;

  wire   [8:1] carry;

  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  XOR2X1 U1 ( .A(B[8]), .B(carry[8]), .Y(SUM[8]) );
  XOR2X1 U2 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
  AND2X1 U3 ( .A(A[0]), .B(B[0]), .Y(carry[1]) );
endmodule


module dacmux_a0_DW01_add_13 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;

  wire   [8:1] carry;

  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  XOR2X1 U1 ( .A(B[8]), .B(carry[8]), .Y(SUM[8]) );
  XOR2X1 U2 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
  AND2X1 U3 ( .A(A[0]), .B(B[0]), .Y(carry[1]) );
endmodule


module dacmux_a0_DW01_add_12 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;

  wire   [8:1] carry;

  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  XOR2X1 U1 ( .A(B[8]), .B(carry[8]), .Y(SUM[8]) );
  AND2X1 U2 ( .A(A[0]), .B(B[0]), .Y(carry[1]) );
  XOR2XL U3 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
endmodule


module dacmux_a0_DW01_add_11 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;

  wire   [8:1] carry;

  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  XOR2X1 U1 ( .A(B[8]), .B(carry[8]), .Y(SUM[8]) );
  XOR2X1 U2 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
  AND2X1 U3 ( .A(A[0]), .B(B[0]), .Y(carry[1]) );
endmodule


module dacmux_a0_DW01_add_10 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;

  wire   [8:1] carry;

  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  XOR2X1 U1 ( .A(B[8]), .B(carry[8]), .Y(SUM[8]) );
  XOR2X1 U2 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
  AND2X1 U3 ( .A(A[0]), .B(B[0]), .Y(carry[1]) );
endmodule


module dacmux_a0_DW01_add_9 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;

  wire   [8:1] carry;

  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  XOR2X1 U1 ( .A(B[8]), .B(carry[8]), .Y(SUM[8]) );
  AND2X1 U2 ( .A(A[0]), .B(B[0]), .Y(carry[1]) );
  XOR2XL U3 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
endmodule


module dacmux_a0_DW01_add_8 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;

  wire   [8:1] carry;

  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  XOR2X1 U1 ( .A(B[8]), .B(carry[8]), .Y(SUM[8]) );
  AND2X1 U2 ( .A(A[0]), .B(B[0]), .Y(carry[1]) );
  XOR2XL U3 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
endmodule


module dacmux_a0_DW01_add_7 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;

  wire   [8:1] carry;

  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  XOR2X1 U1 ( .A(B[8]), .B(carry[8]), .Y(SUM[8]) );
  AND2X1 U2 ( .A(A[0]), .B(B[0]), .Y(carry[1]) );
  XOR2XL U3 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
endmodule


module dacmux_a0_DW01_add_6 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;

  wire   [8:1] carry;

  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  XOR2X1 U1 ( .A(B[8]), .B(carry[8]), .Y(SUM[8]) );
  AND2X1 U2 ( .A(A[0]), .B(B[0]), .Y(carry[1]) );
  XOR2XL U3 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
endmodule


module dacmux_a0_DW01_add_5 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;

  wire   [8:1] carry;

  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  XOR2X1 U1 ( .A(B[8]), .B(carry[8]), .Y(SUM[8]) );
  AND2X1 U2 ( .A(A[0]), .B(B[0]), .Y(carry[1]) );
  XOR2XL U3 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
endmodule


module dacmux_a0_DW01_add_4 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;

  wire   [8:1] carry;

  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  XOR2X1 U1 ( .A(B[8]), .B(carry[8]), .Y(SUM[8]) );
  AND2X1 U2 ( .A(A[0]), .B(B[0]), .Y(carry[1]) );
  XOR2XL U3 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
endmodule


module dacmux_a0_DW01_add_3 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;

  wire   [8:1] carry;

  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  XOR2X1 U1 ( .A(B[8]), .B(carry[8]), .Y(SUM[8]) );
  AND2X1 U2 ( .A(A[0]), .B(B[0]), .Y(carry[1]) );
  XOR2XL U3 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
endmodule


module dacmux_a0_DW01_add_2 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;

  wire   [8:1] carry;

  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  XOR2X1 U1 ( .A(B[8]), .B(carry[8]), .Y(SUM[8]) );
  AND2X1 U2 ( .A(A[0]), .B(B[0]), .Y(carry[1]) );
  XOR2XL U3 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
endmodule


module dacmux_a0_DW01_add_1 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;

  wire   [8:1] carry;

  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  XOR2X1 U1 ( .A(B[8]), .B(carry[8]), .Y(SUM[8]) );
  AND2X1 U2 ( .A(A[0]), .B(B[0]), .Y(carry[1]) );
  XOR2XL U3 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
endmodule


module dacmux_a0_DW01_add_0 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;

  wire   [8:1] carry;

  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  XOR2X1 U1 ( .A(B[8]), .B(carry[8]), .Y(SUM[8]) );
  AND2X1 U2 ( .A(A[0]), .B(B[0]), .Y(carry[1]) );
  XOR2XL U3 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
endmodule


module glreg_WIDTH2_0 ( clk, arstz, we, wdat, rdat );
  input [1:0] wdat;
  output [1:0] rdat;
  input clk, arstz, we;
  wire   n1, n4, n5;

  DFFRQX1 mem_reg_1_ ( .D(n4), .C(clk), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_0_ ( .D(n5), .C(clk), .XR(arstz), .Q(rdat[0]) );
  INVX1 U2 ( .A(we), .Y(n1) );
  AO22XL U3 ( .A(we), .B(wdat[0]), .C(rdat[0]), .D(n1), .Y(n5) );
  AO22XL U4 ( .A(wdat[1]), .B(we), .C(rdat[1]), .D(n1), .Y(n4) );
endmodule


module glreg_WIDTH2_1 ( clk, arstz, we, wdat, rdat );
  input [1:0] wdat;
  output [1:0] rdat;
  input clk, arstz, we;
  wire   n8, n1, n5, n6, n7;

  DFFRQX1 mem_reg_0_ ( .D(n7), .C(clk), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_1_ ( .D(n6), .C(clk), .XR(arstz), .Q(n8) );
  INVXL U2 ( .A(n8), .Y(n1) );
  INVXL U3 ( .A(n1), .Y(rdat[1]) );
  INVXL U4 ( .A(we), .Y(n5) );
  AO22XL U5 ( .A(we), .B(wdat[0]), .C(rdat[0]), .D(n5), .Y(n7) );
  AO22XL U6 ( .A(wdat[1]), .B(we), .C(n8), .D(n5), .Y(n6) );
endmodule


module glreg_a0_25 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net9677;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_25 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9677), .TE(1'b0) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net9677), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net9677), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net9677), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net9677), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net9677), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net9677), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net9677), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net9677), .XR(arstz), .Q(rdat[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_25 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_26 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net9695;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_26 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9695), .TE(1'b0) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net9695), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net9695), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net9695), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net9695), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net9695), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net9695), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net9695), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net9695), .XR(arstz), .Q(rdat[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_26 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_27 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net9713;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_27 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9713), .TE(1'b0) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net9713), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net9713), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net9713), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net9713), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net9713), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net9713), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net9713), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net9713), .XR(arstz), .Q(rdat[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_27 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_28 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net9731;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_28 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9731), .TE(1'b0) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net9731), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net9731), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net9731), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net9731), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net9731), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net9731), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net9731), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net9731), .XR(arstz), .Q(rdat[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_28 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glsta_a0_1 ( clk, arstz, rst0, set2, clr1, rdat, irq );
  input [7:0] set2;
  input [7:0] clr1;
  output [7:0] rdat;
  output [7:0] irq;
  input clk, arstz, rst0;
  wire   upd_r, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22;
  wire   [7:0] wd_r;

  glreg_WIDTH8_1 u0 ( .clk(clk), .arstz(arstz), .we(upd_r), .wdat(wd_r), 
        .rdat(rdat) );
  INVX1 U2 ( .A(set2[4]), .Y(n14) );
  INVX1 U3 ( .A(set2[5]), .Y(n9) );
  NAND31X1 U4 ( .C(set2[5]), .A(n8), .B(n7), .Y(n1) );
  NOR8XL U5 ( .A(clr1[3]), .B(clr1[2]), .C(clr1[1]), .D(clr1[0]), .E(clr1[7]), 
        .F(clr1[6]), .G(clr1[5]), .H(clr1[4]), .Y(n4) );
  INVX1 U6 ( .A(set2[6]), .Y(n8) );
  INVX1 U7 ( .A(set2[7]), .Y(n7) );
  INVX1 U8 ( .A(set2[0]), .Y(n10) );
  INVX1 U9 ( .A(set2[2]), .Y(n12) );
  INVX1 U10 ( .A(set2[1]), .Y(n11) );
  INVX1 U11 ( .A(set2[3]), .Y(n13) );
  NAND42X1 U12 ( .C(n6), .D(n5), .A(n4), .B(n3), .Y(upd_r) );
  NOR32XL U13 ( .B(n14), .C(n2), .A(n1), .Y(n3) );
  NAND21X1 U14 ( .B(set2[3]), .A(n12), .Y(n6) );
  NAND21X1 U15 ( .B(set2[1]), .A(n10), .Y(n5) );
  AOI211X1 U16 ( .C(n8), .D(n16), .A(rst0), .B(clr1[6]), .Y(wd_r[6]) );
  INVX1 U17 ( .A(rdat[6]), .Y(n16) );
  AOI211X1 U18 ( .C(n7), .D(n15), .A(rst0), .B(clr1[7]), .Y(wd_r[7]) );
  INVX1 U19 ( .A(rdat[7]), .Y(n15) );
  AOI211X1 U20 ( .C(n11), .D(n21), .A(rst0), .B(clr1[1]), .Y(wd_r[1]) );
  INVX1 U21 ( .A(rdat[1]), .Y(n21) );
  AOI211X1 U22 ( .C(n12), .D(n20), .A(rst0), .B(clr1[2]), .Y(wd_r[2]) );
  INVX1 U23 ( .A(rdat[2]), .Y(n20) );
  AOI211X1 U24 ( .C(n14), .D(n18), .A(rst0), .B(clr1[4]), .Y(wd_r[4]) );
  INVX1 U25 ( .A(rdat[4]), .Y(n18) );
  AOI211X1 U26 ( .C(n9), .D(n17), .A(rst0), .B(clr1[5]), .Y(wd_r[5]) );
  INVX1 U27 ( .A(rdat[5]), .Y(n17) );
  AOI211X1 U28 ( .C(n10), .D(n22), .A(rst0), .B(clr1[0]), .Y(wd_r[0]) );
  INVX1 U29 ( .A(rdat[0]), .Y(n22) );
  AOI211X1 U30 ( .C(n13), .D(n19), .A(rst0), .B(clr1[3]), .Y(wd_r[3]) );
  INVX1 U31 ( .A(rdat[3]), .Y(n19) );
  NOR2X1 U32 ( .A(rdat[3]), .B(n13), .Y(irq[3]) );
  NOR2X1 U33 ( .A(rdat[2]), .B(n12), .Y(irq[2]) );
  NOR2X1 U34 ( .A(rdat[1]), .B(n11), .Y(irq[1]) );
  NOR2X1 U35 ( .A(rdat[5]), .B(n9), .Y(irq[5]) );
  NOR2X1 U36 ( .A(rdat[0]), .B(n10), .Y(irq[0]) );
  NOR2X1 U37 ( .A(rdat[4]), .B(n14), .Y(irq[4]) );
  NOR2X1 U38 ( .A(rdat[6]), .B(n8), .Y(irq[6]) );
  NOR2X1 U39 ( .A(rdat[7]), .B(n7), .Y(irq[7]) );
  INVX1 U40 ( .A(rst0), .Y(n2) );
endmodule


module glreg_WIDTH8_1 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net9749;

  SNPS_CLOCK_GATE_HIGH_glreg_WIDTH8_1 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9749), .TE(1'b0) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net9749), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net9749), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net9749), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net9749), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net9749), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net9749), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net9749), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net9749), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_WIDTH8_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_29 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net9767;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_29 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9767), .TE(1'b0) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net9767), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net9767), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net9767), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net9767), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net9767), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net9767), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net9767), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net9767), .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_29 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_30 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net9785;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_30 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9785), .TE(1'b0) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net9785), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net9785), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net9785), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net9785), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net9785), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net9785), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net9785), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net9785), .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_30 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_31 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net9803;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_31 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9803), .TE(1'b0) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net9803), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net9803), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net9803), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net9803), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net9803), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net9803), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net9803), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net9803), .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_31 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_32 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net9821;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_32 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9821), .TE(1'b0) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net9821), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net9821), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net9821), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net9821), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net9821), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net9821), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net9821), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net9821), .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_32 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_33 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net9839;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_33 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9839), .TE(1'b0) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net9839), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net9839), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net9839), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net9839), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net9839), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net9839), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net9839), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net9839), .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_33 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_34 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net9857;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_34 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9857), .TE(1'b0) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net9857), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net9857), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net9857), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net9857), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net9857), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net9857), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net9857), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net9857), .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_34 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_35 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net9875;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_35 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9875), .TE(1'b0) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net9875), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net9875), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net9875), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net9875), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net9875), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net9875), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net9875), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net9875), .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_35 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_36 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net9893;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_36 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9893), .TE(1'b0) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net9893), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net9893), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net9893), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net9893), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net9893), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net9893), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net9893), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net9893), .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_36 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_37 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net9911;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_37 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9911), .TE(1'b0) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net9911), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net9911), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net9911), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net9911), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net9911), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net9911), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net9911), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net9911), .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_37 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_38 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net9929;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_38 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9929), .TE(1'b0) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net9929), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net9929), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net9929), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net9929), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net9929), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net9929), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net9929), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net9929), .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_38 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_39 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net9947;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_39 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9947), .TE(1'b0) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net9947), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net9947), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net9947), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net9947), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net9947), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net9947), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net9947), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net9947), .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_39 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_40 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net9965;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_40 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9965), .TE(1'b0) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net9965), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net9965), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net9965), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net9965), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net9965), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net9965), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net9965), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net9965), .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_40 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_41 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net9983;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_41 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net9983), .TE(1'b0) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net9983), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net9983), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net9983), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net9983), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net9983), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net9983), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net9983), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net9983), .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_41 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_42 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net10001;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_42 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10001), .TE(1'b0) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net10001), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net10001), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net10001), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net10001), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net10001), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net10001), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net10001), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net10001), .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_42 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_43 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net10019;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_43 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10019), .TE(1'b0) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net10019), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net10019), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net10019), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net10019), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net10019), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net10019), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net10019), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net10019), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_43 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_44 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net10037;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_44 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10037), .TE(1'b0) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net10037), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net10037), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net10037), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net10037), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net10037), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net10037), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net10037), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net10037), .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_44 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_45 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net10055;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_45 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10055), .TE(1'b0) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net10055), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net10055), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net10055), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net10055), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net10055), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net10055), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net10055), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net10055), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_45 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_46 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net10073;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_46 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10073), .TE(1'b0) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net10073), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net10073), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net10073), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net10073), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net10073), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net10073), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net10073), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net10073), .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_46 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_WIDTH6_2 ( clk, arstz, we, wdat, rdat );
  input [5:0] wdat;
  output [5:0] rdat;
  input clk, arstz, we;
  wire   net10091;

  SNPS_CLOCK_GATE_HIGH_glreg_WIDTH6_2 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10091), .TE(1'b0) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net10091), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net10091), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net10091), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net10091), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net10091), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net10091), .XR(arstz), .Q(rdat[3]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_WIDTH6_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_47 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net10109;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_47 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10109), .TE(1'b0) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net10109), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net10109), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net10109), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net10109), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net10109), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net10109), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net10109), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net10109), .XR(arstz), .Q(rdat[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_47 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_48 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net10127;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_48 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10127), .TE(1'b0) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net10127), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net10127), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net10127), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net10127), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net10127), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net10127), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net10127), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net10127), .XR(arstz), .Q(rdat[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_48 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_WIDTH7_1 ( clk, arstz, we, wdat, rdat );
  input [6:0] wdat;
  output [6:0] rdat;
  input clk, arstz, we;
  wire   net10145;

  SNPS_CLOCK_GATE_HIGH_glreg_WIDTH7_1 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10145), .TE(1'b0) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net10145), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net10145), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net10145), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net10145), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net10145), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net10145), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net10145), .XR(arstz), .Q(rdat[6]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_WIDTH7_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module shmux_00000005_00000012_00000012 ( ps_sample, ps_md4ch, r_comp_swtch, 
        r_semi, r_loop, r_dac_en, wr_dacv, busy, sh_hold, stop, semi_start, 
        auto_start, mxcyc_done, sampl_begn, sampl_done, app_dacis, pos_dacis, 
        cs_ptr, ps_ptr, clk, srstz );
  input [17:0] r_dac_en;
  input [17:0] wr_dacv;
  output [17:0] app_dacis;
  output [17:0] pos_dacis;
  output [4:0] cs_ptr;
  output [4:0] ps_ptr;
  input ps_sample, ps_md4ch, r_comp_swtch, r_semi, r_loop, stop, semi_start,
         auto_start, mxcyc_done, sampl_begn, sampl_done, clk, srstz;
  output busy, sh_hold;
  wire   n760, cs_mux_5_, N956, N957, N958, N959, N960, N961, N962, N963, N964,
         N965, N966, N967, N968, N969, N970, N971, N972, N973, N1002, N1003,
         N1004, N1005, N1006, N1007, N1008, N1009, N1010, N1011, N1012, N1013,
         N1014, N1015, N1016, N1017, N1018, N1019, N1020, N1030, N1031, N1032,
         N1033, N1034, N1035, N1172, N1173, N1174, N1175, N1176, N1181, N1182,
         N1183, N1184, N1185, N1215, N1217, N1222, N1223, N1224, N1225, N1226,
         N1254, N1255, N1256, N1257, N1258, N1263, N1264, N1265, N1266, N1267,
         N1296, N1297, N1298, N1299, N1304, N1305, N1306, N1307, N1308, N1336,
         N1337, N1338, N1339, N1340, N1345, N1346, N1347, N1348, N1349, N1379,
         N1380, N1381, N1386, N1387, N1388, N1389, N1390, N1418, N1419, N1420,
         N1421, N1422, N1427, N1428, N1429, N1430, N1431, N1460, N1461, N1462,
         N1463, N1464, N1472, N1500, N1501, N1502, N1503, N1504, N1505, N1509,
         N1513, N1542, N1544, N1545, N1546, N1550, N1552, N1582, N1583, N1584,
         N1585, N1586, N1591, N1592, N1593, N1594, N1595, N1624, N1625, N1626,
         N1627, N1628, N1636, N1664, N1665, N1666, N1667, N1668, N1669, N1673,
         N1677, N1705, N1707, N1708, N1709, N1714, N1715, N1716, N1717, N1718,
         N1750, N1755, N1756, N1795, N1796, N1797, N1837, N1838, net10163,
         net10169, n284, n285, n286, n287, n288, n289, n301, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n322,
         n334, n338, n339, n340, n341, n342, n343, n358, n359, n360, n361,
         n375, n376, n377, n378, n397, n398, n399, n400, n419, n420, n421,
         n422, n423, n424, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n660, add_394_carry_2_,
         add_394_carry_3_, add_394_carry_4_, add_394_I3_carry_2_,
         add_394_I3_carry_3_, add_394_I3_carry_4_, add_394_I5_carry_2_,
         add_394_I5_carry_3_, add_394_I5_carry_4_, add_394_I6_carry_4_,
         add_394_I7_carry_2_, add_394_I7_carry_3_, add_394_I7_carry_4_,
         add_394_I9_carry_2_, add_394_I9_carry_3_, add_394_I9_carry_4_,
         add_394_I11_carry_2_, add_394_I11_carry_3_, add_394_I11_carry_4_,
         add_394_I13_carry_2_, add_394_I13_carry_3_, add_394_I13_carry_4_,
         add_394_I14_carry_4_, add_394_I15_carry_2_, add_394_I15_carry_3_,
         add_394_I15_carry_4_, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n76, n77, n78, n79, n80, n81, n83, n84,
         n85, n86, n87, n89, n90, n91, n92, n93, n95, n96, n97, n98, n99, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n302, n303, n317, n318, n319,
         n320, n321, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n335, n336, n337, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n425, n608, n609, n610, n611, n612, n613, n614, n625,
         n626, n627, n628, n639, n640, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759;
  wire   [17:0] neg_dacis;
  wire   [5:2] sub_395_S2_aco_carry;
  wire   [5:2] sub_395_S2_I2_aco_carry;
  wire   [5:2] sub_395_S2_I3_aco_carry;
  wire   [5:2] sub_395_S2_I4_aco_carry;
  wire   [4:3] add_394_I4_carry;
  wire   [5:2] sub_395_S2_I5_aco_carry;
  wire   [5:2] sub_395_S2_I6_aco_carry;
  wire   [5:2] sub_395_S2_I7_aco_carry;
  wire   [5:2] sub_395_S2_I8_aco_carry;
  wire   [4:3] add_394_I8_carry;
  wire   [5:2] sub_395_S2_I9_aco_carry;
  wire   [5:2] sub_395_S2_I10_aco_carry;
  wire   [5:2] sub_395_S2_I11_aco_carry;
  wire   [5:2] sub_395_S2_I12_aco_carry;
  wire   [4:3] add_394_I12_carry;
  wire   [5:2] sub_395_S2_I13_aco_carry;
  wire   [5:2] sub_395_S2_I14_aco_carry;
  wire   [4:3] add_394_I16_carry;

  SNPS_CLOCK_GATE_HIGH_shmux_00000005_00000012_00000012_0 clk_gate_r_dacis_reg ( 
        .CLK(clk), .EN(N1002), .ENCLK(net10163), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_shmux_00000005_00000012_00000012_1 clk_gate_cs_mux_reg ( 
        .CLK(clk), .EN(N1030), .ENCLK(net10169), .TE(1'b0) );
  FAD1X1 sub_395_S2_aco_U2_4 ( .A(N1175), .B(n55), .CI(sub_395_S2_aco_carry[4]), .CO(sub_395_S2_aco_carry[5]), .SO(N1184) );
  FAD1X1 sub_395_S2_I2_aco_U2_4 ( .A(n103), .B(n71), .CI(
        sub_395_S2_I2_aco_carry[4]), .CO(sub_395_S2_I2_aco_carry[5]), .SO(
        N1225) );
  FAD1X1 sub_395_S2_I3_aco_U2_4 ( .A(N1257), .B(n56), .CI(
        sub_395_S2_I3_aco_carry[4]), .CO(sub_395_S2_I3_aco_carry[5]), .SO(
        N1266) );
  FAD1X1 sub_395_S2_I4_aco_U2_4 ( .A(N1298), .B(n67), .CI(
        sub_395_S2_I4_aco_carry[4]), .CO(sub_395_S2_I4_aco_carry[5]), .SO(
        N1307) );
  FAD1X1 sub_395_S2_I5_aco_U2_4 ( .A(N1339), .B(n54), .CI(
        sub_395_S2_I5_aco_carry[4]), .CO(sub_395_S2_I5_aco_carry[5]), .SO(
        N1348) );
  FAD1X1 sub_395_S2_I6_aco_U2_4 ( .A(N1380), .B(n68), .CI(
        sub_395_S2_I6_aco_carry[4]), .CO(sub_395_S2_I6_aco_carry[5]), .SO(
        N1389) );
  FAD1X1 sub_395_S2_I7_aco_U2_4 ( .A(N1421), .B(n52), .CI(
        sub_395_S2_I7_aco_carry[4]), .CO(sub_395_S2_I7_aco_carry[5]), .SO(
        N1430) );
  FAD1X1 sub_395_S2_I11_aco_U2_4 ( .A(N1585), .B(n53), .CI(
        sub_395_S2_I11_aco_carry[4]), .CO(sub_395_S2_I11_aco_carry[5]), .SO(
        N1594) );
  FAD1X1 sub_395_S2_I14_aco_U2_4 ( .A(N1708), .B(n66), .CI(
        sub_395_S2_I14_aco_carry[4]), .CO(sub_395_S2_I14_aco_carry[5]), .SO(
        N1717) );
  DFFQX1 cs_mux_reg_1_ ( .D(N1032), .C(net10169), .Q(N1705) );
  DFFQX1 cs_mux_reg_2_ ( .D(N1033), .C(net10169), .Q(N1542) );
  DFFQX1 cs_mux_reg_3_ ( .D(N1034), .C(net10169), .Q(N1215) );
  DFFQX1 cs_mux_reg_4_ ( .D(N1035), .C(net10169), .Q(N1217) );
  DFFQX1 cs_mux_reg_0_ ( .D(N1031), .C(net10169), .Q(N1795) );
  DFFQX1 r_dacis_reg_16_ ( .D(N1019), .C(net10163), .Q(pos_dacis[16]) );
  DFFQX1 r_dacis_reg_11_ ( .D(N1014), .C(net10163), .Q(pos_dacis[11]) );
  DFFQX1 r_dacis_reg_13_ ( .D(N1016), .C(net10163), .Q(pos_dacis[13]) );
  DFFQX1 r_dacis_reg_10_ ( .D(N1013), .C(net10163), .Q(pos_dacis[10]) );
  DFFQX1 r_dacis_reg_17_ ( .D(N1020), .C(net10163), .Q(pos_dacis[17]) );
  DFFQX1 r_dacis_reg_15_ ( .D(N1018), .C(net10163), .Q(pos_dacis[15]) );
  DFFQX1 r_dacis_reg_12_ ( .D(N1015), .C(net10163), .Q(pos_dacis[12]) );
  DFFQX1 r_dacis_reg_14_ ( .D(N1017), .C(net10163), .Q(pos_dacis[14]) );
  DFFQX1 r_dacis_reg_9_ ( .D(N1012), .C(net10163), .Q(pos_dacis[9]) );
  DFFQX1 r_dacis_reg_8_ ( .D(N1011), .C(net10163), .Q(pos_dacis[8]) );
  DFFNQX1 neg_dacis_reg_0_ ( .D(N956), .XC(clk), .Q(neg_dacis[0]) );
  DFFNQX1 neg_dacis_reg_1_ ( .D(N957), .XC(clk), .Q(neg_dacis[1]) );
  DFFNQX1 neg_dacis_reg_2_ ( .D(N958), .XC(clk), .Q(neg_dacis[2]) );
  DFFNQX1 neg_dacis_reg_3_ ( .D(N959), .XC(clk), .Q(neg_dacis[3]) );
  DFFNQX1 neg_dacis_reg_4_ ( .D(N960), .XC(clk), .Q(neg_dacis[4]) );
  DFFNQX1 neg_dacis_reg_5_ ( .D(N961), .XC(clk), .Q(neg_dacis[5]) );
  DFFNQX1 neg_dacis_reg_6_ ( .D(N962), .XC(clk), .Q(neg_dacis[6]) );
  DFFNQX1 neg_dacis_reg_7_ ( .D(N963), .XC(clk), .Q(neg_dacis[7]) );
  DFFNQX1 neg_dacis_reg_8_ ( .D(N964), .XC(clk), .Q(neg_dacis[8]) );
  DFFNQX1 neg_dacis_reg_9_ ( .D(N965), .XC(clk), .Q(neg_dacis[9]) );
  DFFNQX1 neg_dacis_reg_10_ ( .D(N966), .XC(clk), .Q(neg_dacis[10]) );
  DFFNQX1 neg_dacis_reg_11_ ( .D(N967), .XC(clk), .Q(neg_dacis[11]) );
  DFFNQX1 neg_dacis_reg_12_ ( .D(N968), .XC(clk), .Q(neg_dacis[12]) );
  DFFNQX1 neg_dacis_reg_13_ ( .D(N969), .XC(clk), .Q(neg_dacis[13]) );
  DFFNQX1 neg_dacis_reg_14_ ( .D(N970), .XC(clk), .Q(neg_dacis[14]) );
  DFFNQX1 neg_dacis_reg_15_ ( .D(N971), .XC(clk), .Q(neg_dacis[15]) );
  DFFNQX1 neg_dacis_reg_16_ ( .D(N972), .XC(clk), .Q(neg_dacis[16]) );
  DFFNQX1 neg_dacis_reg_17_ ( .D(N973), .XC(clk), .Q(neg_dacis[17]) );
  DFFQX1 cs_mux_reg_5_ ( .D(n660), .C(clk), .Q(cs_mux_5_) );
  DFFQX1 r_dacis_reg_7_ ( .D(N1010), .C(net10163), .Q(pos_dacis[7]) );
  DFFQX1 r_dacis_reg_6_ ( .D(N1009), .C(net10163), .Q(pos_dacis[6]) );
  DFFQX1 r_dacis_reg_5_ ( .D(N1008), .C(net10163), .Q(pos_dacis[5]) );
  DFFQX1 r_dacis_reg_4_ ( .D(N1007), .C(net10163), .Q(pos_dacis[4]) );
  DFFQX1 r_dacis_reg_2_ ( .D(N1005), .C(net10163), .Q(pos_dacis[2]) );
  DFFQX1 r_dacis_reg_3_ ( .D(N1006), .C(net10163), .Q(pos_dacis[3]) );
  DFFQX1 r_dacis_reg_1_ ( .D(N1004), .C(net10163), .Q(pos_dacis[1]) );
  DFFQX1 r_dacis_reg_0_ ( .D(N1003), .C(net10163), .Q(pos_dacis[0]) );
  NAND32X1 U3 ( .B(n69), .C(n188), .A(n112), .Y(n111) );
  INVX1 U4 ( .A(n407), .Y(n167) );
  GEN2XL U5 ( .D(n232), .E(n91), .C(n231), .B(n235), .A(n201), .Y(n175) );
  GEN3XL U6 ( .F(n264), .G(n263), .E(n262), .D(n261), .C(n260), .B(n259), .A(
        n258), .Y(n265) );
  OA2222XL U7 ( .A(n164), .B(n273), .C(n163), .D(n370), .E(n162), .F(n269), 
        .G(n161), .H(n369), .Y(n169) );
  AOI31X1 U8 ( .A(n339), .B(n340), .C(n338), .D(n281), .Y(n241) );
  NAND42X1 U9 ( .C(n229), .D(n228), .A(n227), .B(n226), .Y(ps_ptr[3]) );
  OA222X1 U10 ( .A(n3), .B(n271), .C(n62), .D(n383), .E(n57), .F(n274), .Y(
        n226) );
  NAND43X1 U11 ( .B(n216), .C(n215), .D(n65), .A(n214), .Y(ps_ptr[1]) );
  AND4X1 U12 ( .A(n73), .B(n207), .C(n206), .D(n32), .Y(n216) );
  OAI222XL U13 ( .A(n665), .B(n271), .C(n673), .D(n383), .E(n669), .F(n274), 
        .Y(n1) );
  MUX2IX1 U14 ( .D0(N1217), .D1(ps_ptr[4]), .S(ps_sample), .Y(n2) );
  OA22X1 U15 ( .A(n148), .B(n147), .C(n146), .D(n145), .Y(n3) );
  INVX1 U16 ( .A(n245), .Y(n4) );
  INVX1 U17 ( .A(r_dac_en[16]), .Y(n5) );
  INVX1 U18 ( .A(n5), .Y(n6) );
  INVX1 U19 ( .A(n5), .Y(n7) );
  INVX1 U20 ( .A(r_dac_en[0]), .Y(n8) );
  INVX1 U21 ( .A(n8), .Y(n9) );
  INVX1 U22 ( .A(n8), .Y(n10) );
  INVX1 U23 ( .A(r_dac_en[3]), .Y(n11) );
  INVX1 U24 ( .A(n11), .Y(n12) );
  INVX1 U25 ( .A(n11), .Y(n13) );
  INVX1 U26 ( .A(r_dac_en[9]), .Y(n14) );
  INVX1 U27 ( .A(n14), .Y(n15) );
  INVX1 U28 ( .A(n14), .Y(n16) );
  INVX1 U29 ( .A(r_dac_en[10]), .Y(n17) );
  INVX1 U30 ( .A(n17), .Y(n18) );
  INVX1 U31 ( .A(n17), .Y(n19) );
  INVX1 U32 ( .A(r_dac_en[11]), .Y(n20) );
  INVX1 U33 ( .A(n20), .Y(n21) );
  INVX1 U34 ( .A(n20), .Y(n22) );
  INVX1 U35 ( .A(r_dac_en[12]), .Y(n23) );
  INVX1 U36 ( .A(n23), .Y(n24) );
  INVX1 U37 ( .A(n23), .Y(n25) );
  INVX1 U38 ( .A(r_dac_en[13]), .Y(n26) );
  INVX1 U39 ( .A(n26), .Y(n27) );
  INVX1 U40 ( .A(n26), .Y(n28) );
  INVX1 U41 ( .A(r_dac_en[15]), .Y(n29) );
  INVX1 U42 ( .A(n29), .Y(n30) );
  INVX1 U43 ( .A(n29), .Y(n31) );
  INVX1 U44 ( .A(r_dac_en[1]), .Y(n32) );
  INVX1 U45 ( .A(n32), .Y(n33) );
  INVX1 U46 ( .A(n32), .Y(n34) );
  INVX1 U47 ( .A(r_dac_en[2]), .Y(n35) );
  INVX1 U48 ( .A(n35), .Y(n36) );
  INVX1 U49 ( .A(n35), .Y(n37) );
  INVX1 U50 ( .A(r_dac_en[8]), .Y(n38) );
  INVX1 U51 ( .A(n38), .Y(n39) );
  INVX1 U52 ( .A(n38), .Y(n40) );
  INVX1 U53 ( .A(r_dac_en[14]), .Y(n41) );
  INVX1 U54 ( .A(n41), .Y(n42) );
  INVX1 U55 ( .A(n41), .Y(n43) );
  INVX1 U56 ( .A(r_dac_en[5]), .Y(n44) );
  INVX1 U57 ( .A(r_dac_en[4]), .Y(n45) );
  INVX1 U58 ( .A(r_dac_en[7]), .Y(n46) );
  INVX1 U59 ( .A(r_dac_en[6]), .Y(n47) );
  NAND2X1 U60 ( .A(sampl_done), .B(srstz), .Y(n48) );
  OA222X1 U61 ( .A(n668), .B(n271), .C(n676), .D(n383), .E(n672), .F(n274), 
        .Y(n214) );
  NAND32X1 U62 ( .B(n154), .C(n179), .A(n180), .Y(n383) );
  OR4X2 U63 ( .A(n242), .B(n241), .C(n59), .D(n1), .Y(ps_ptr[4]) );
  NAND2X1 U64 ( .A(n179), .B(n180), .Y(n274) );
  INVXL U65 ( .A(n383), .Y(n384) );
  NOR43XL U66 ( .B(n249), .C(n248), .D(n41), .A(n50), .Y(n197) );
  INVX1 U67 ( .A(n353), .Y(n356) );
  GEN2XL U68 ( .D(n257), .E(n256), .C(n255), .B(n254), .A(n253), .Y(n263) );
  AND2XL U69 ( .A(n364), .B(n366), .Y(N1004) );
  AND2XL U70 ( .A(n362), .B(n366), .Y(N1006) );
  AND2XL U71 ( .A(n363), .B(n366), .Y(N1005) );
  AND2XL U72 ( .A(n354), .B(n362), .Y(N1014) );
  AND2XL U73 ( .A(n391), .B(ps_ptr[2]), .Y(N1033) );
  AO21XL U74 ( .B(n169), .C(n49), .A(n275), .Y(n170) );
  OA222X1 U75 ( .A(n272), .B(n168), .C(n167), .D(n268), .E(n334), .F(n166), 
        .Y(n49) );
  AND3XL U76 ( .A(n271), .B(n383), .C(n270), .Y(n278) );
  NAND32XL U77 ( .B(n352), .C(n346), .A(n2), .Y(n330) );
  INVXL U78 ( .A(n295), .Y(n299) );
  INVXL U79 ( .A(n351), .Y(n346) );
  NAND21XL U80 ( .B(n2), .A(n346), .Y(n326) );
  AND3XL U81 ( .A(n367), .B(n352), .C(n329), .Y(N1019) );
  AND3XL U82 ( .A(n364), .B(n352), .C(n329), .Y(N1020) );
  OAI21X1 U83 ( .B(n87), .C(n221), .A(n29), .Y(n50) );
  NOR32XL U84 ( .B(n245), .C(n79), .A(wr_dacv[17]), .Y(n246) );
  INVXL U85 ( .A(n231), .Y(n220) );
  OAI211XL U86 ( .C(n98), .D(n221), .A(n220), .B(n235), .Y(n222) );
  INVXL U87 ( .A(n243), .Y(n264) );
  INVXL U88 ( .A(n221), .Y(n232) );
  INVXL U89 ( .A(n253), .Y(n200) );
  INVXL U90 ( .A(n293), .Y(n300) );
  INVXL U91 ( .A(n244), .Y(n257) );
  MUX2XL U92 ( .D0(n77), .D1(ps_ptr[0]), .S(ps_sample), .Y(n344) );
  NAND32XL U93 ( .B(n351), .C(n347), .A(n2), .Y(n357) );
  NAND32XL U94 ( .B(n346), .C(n347), .A(n2), .Y(n348) );
  AND3XL U95 ( .A(n356), .B(n367), .C(n365), .Y(N1007) );
  AND3XL U96 ( .A(n356), .B(n364), .C(n365), .Y(N1008) );
  AND2XL U97 ( .A(n391), .B(ps_ptr[0]), .Y(N1031) );
  NOR3X2 U98 ( .A(wr_dacv[0]), .B(n178), .C(n10), .Y(n73) );
  NAND41XL U99 ( .D(n36), .A(n51), .B(n266), .C(n205), .Y(n206) );
  OAI21X1 U100 ( .B(n204), .C(n203), .A(n217), .Y(n51) );
  INVX1 U101 ( .A(srstz), .Y(n105) );
  INVX1 U102 ( .A(n566), .Y(n693) );
  INVX1 U103 ( .A(n565), .Y(n692) );
  INVX1 U104 ( .A(n494), .Y(n710) );
  INVX1 U105 ( .A(n493), .Y(n709) );
  INVX1 U106 ( .A(n469), .Y(n719) );
  INVX1 U107 ( .A(n470), .Y(n720) );
  INVX1 U108 ( .A(n518), .Y(n730) );
  INVX1 U109 ( .A(n446), .Y(n740) );
  INVX1 U110 ( .A(n517), .Y(n729) );
  INVX1 U111 ( .A(n445), .Y(n739) );
  INVX1 U112 ( .A(n542), .Y(n701) );
  INVX1 U113 ( .A(n603), .Y(n685) );
  INVX1 U114 ( .A(n541), .Y(n700) );
  INVX1 U115 ( .A(n602), .Y(n684) );
  INVX1 U116 ( .A(n145), .Y(n148) );
  INVX1 U117 ( .A(n619), .Y(n674) );
  INVX1 U118 ( .A(n646), .Y(n667) );
  INVX1 U119 ( .A(n645), .Y(n666) );
  INVX1 U120 ( .A(wr_dacv[15]), .Y(n248) );
  INVX1 U121 ( .A(n110), .Y(n391) );
  NAND32X1 U122 ( .B(n109), .C(n105), .A(n302), .Y(n110) );
  INVX1 U123 ( .A(n283), .Y(n109) );
  AO21X1 U124 ( .B(n105), .C(n302), .A(n391), .Y(N1030) );
  INVX1 U125 ( .A(wr_dacv[2]), .Y(n266) );
  INVX1 U126 ( .A(wr_dacv[1]), .Y(n207) );
  INVX1 U127 ( .A(N1505), .Y(n414) );
  INVX1 U128 ( .A(N1669), .Y(n417) );
  INVX1 U129 ( .A(n392), .Y(n682) );
  NOR2X1 U130 ( .A(n694), .B(N1592), .Y(n563) );
  NOR2X1 U131 ( .A(N1591), .B(N1592), .Y(n564) );
  NOR2X1 U132 ( .A(N1427), .B(N1428), .Y(n492) );
  NOR2X1 U133 ( .A(n711), .B(N1428), .Y(n491) );
  INVX1 U134 ( .A(N1345), .Y(n721) );
  INVX1 U135 ( .A(N1263), .Y(n731) );
  INVX1 U136 ( .A(N1591), .Y(n694) );
  INVX1 U137 ( .A(N1427), .Y(n711) );
  INVX1 U138 ( .A(N1594), .Y(n690) );
  INVX1 U139 ( .A(N1430), .Y(n707) );
  INVX1 U140 ( .A(N1348), .Y(n717) );
  INVX1 U141 ( .A(N1266), .Y(n727) );
  NAND2X1 U142 ( .A(N1592), .B(n694), .Y(n565) );
  NAND2XL U143 ( .A(N1592), .B(N1591), .Y(n566) );
  NAND2XL U144 ( .A(N1428), .B(N1427), .Y(n494) );
  NAND2X1 U145 ( .A(N1428), .B(n711), .Y(n493) );
  NAND2X1 U146 ( .A(N1346), .B(n721), .Y(n469) );
  NOR2X1 U147 ( .A(N1345), .B(N1346), .Y(n468) );
  NOR2X1 U148 ( .A(N1263), .B(N1264), .Y(n516) );
  NOR2X1 U149 ( .A(N1181), .B(N1182), .Y(n444) );
  NOR2X1 U150 ( .A(n721), .B(N1346), .Y(n467) );
  NOR2X1 U151 ( .A(n731), .B(N1264), .Y(n515) );
  NOR2X1 U152 ( .A(n741), .B(N1182), .Y(n443) );
  NOR2X1 U153 ( .A(n211), .B(n407), .Y(n600) );
  NOR2X1 U154 ( .A(N1673), .B(n407), .Y(n601) );
  INVX1 U155 ( .A(N1181), .Y(n741) );
  INVX1 U156 ( .A(N1593), .Y(n691) );
  INVX1 U157 ( .A(N1306), .Y(n723) );
  INVX1 U158 ( .A(N1429), .Y(n708) );
  INVX1 U159 ( .A(N1184), .Y(n737) );
  INVX1 U160 ( .A(n211), .Y(N1673) );
  INVX1 U161 ( .A(n208), .Y(N1509) );
  NAND2XL U162 ( .A(N1346), .B(N1345), .Y(n470) );
  NAND2XL U163 ( .A(N1264), .B(N1263), .Y(n518) );
  NAND2XL U164 ( .A(N1182), .B(N1181), .Y(n446) );
  NAND2X1 U165 ( .A(N1264), .B(n731), .Y(n517) );
  NAND2X1 U166 ( .A(N1182), .B(n741), .Y(n445) );
  NAND2X1 U167 ( .A(n411), .B(n208), .Y(n541) );
  NAND2X1 U168 ( .A(n407), .B(n211), .Y(n602) );
  NAND2X1 U169 ( .A(n411), .B(N1509), .Y(n542) );
  NAND2X1 U170 ( .A(n407), .B(N1673), .Y(n603) );
  INVX1 U171 ( .A(n401), .Y(n683) );
  NOR2X1 U172 ( .A(n208), .B(n411), .Y(n539) );
  NOR2X1 U173 ( .A(N1509), .B(n411), .Y(n540) );
  INVX1 U174 ( .A(n123), .Y(n187) );
  INVX1 U175 ( .A(n133), .Y(n121) );
  INVX1 U176 ( .A(n505), .Y(n724) );
  INVX1 U177 ( .A(n578), .Y(n688) );
  INVX1 U178 ( .A(n577), .Y(n687) );
  NAND21X1 U179 ( .B(n132), .A(n191), .Y(n145) );
  INVX1 U180 ( .A(N1837), .Y(n668) );
  NAND2X1 U181 ( .A(N1756), .B(n676), .Y(n619) );
  INVX1 U182 ( .A(n403), .Y(n686) );
  INVX1 U183 ( .A(n404), .Y(n699) );
  NOR2X1 U184 ( .A(n676), .B(N1756), .Y(n617) );
  NOR2X1 U185 ( .A(n668), .B(N1838), .Y(n643) );
  NOR2X1 U186 ( .A(N1837), .B(N1838), .Y(n644) );
  INVX1 U187 ( .A(n138), .Y(n124) );
  INVX1 U188 ( .A(n530), .Y(n704) );
  INVX1 U189 ( .A(n620), .Y(n675) );
  INVX1 U190 ( .A(n529), .Y(n703) );
  INVX1 U191 ( .A(N1592), .Y(n166) );
  NAND2X1 U192 ( .A(N1838), .B(N1837), .Y(n646) );
  NAND2X1 U193 ( .A(N1838), .B(n668), .Y(n645) );
  INVX1 U194 ( .A(n402), .Y(n702) );
  INVX1 U195 ( .A(n458), .Y(n735) );
  INVX1 U196 ( .A(n457), .Y(n734) );
  INVX1 U197 ( .A(n633), .Y(n670) );
  INVX1 U198 ( .A(n396), .Y(n237) );
  INVX1 U199 ( .A(n411), .Y(n162) );
  INVX1 U200 ( .A(wr_dacv[14]), .Y(n249) );
  INVX3 U201 ( .A(auto_start), .Y(n151) );
  INVXL U202 ( .A(ps_ptr[3]), .Y(n320) );
  AND2X1 U203 ( .A(n345), .B(n362), .Y(N1018) );
  AND2X1 U204 ( .A(n345), .B(n363), .Y(N1017) );
  AND2X1 U205 ( .A(n345), .B(n364), .Y(N1016) );
  AND2X1 U206 ( .A(n345), .B(n367), .Y(N1015) );
  AND2X1 U207 ( .A(n356), .B(n362), .Y(N1010) );
  AND2X1 U208 ( .A(n356), .B(n363), .Y(N1009) );
  INVX1 U209 ( .A(wr_dacv[8]), .Y(n199) );
  INVX1 U210 ( .A(n333), .Y(n337) );
  NAND21X1 U211 ( .B(n332), .A(n331), .Y(n333) );
  NAND32XL U212 ( .B(mxcyc_done), .C(semi_start), .A(n151), .Y(n283) );
  INVX1 U213 ( .A(n350), .Y(n367) );
  INVX1 U214 ( .A(n336), .Y(n362) );
  NAND21X1 U215 ( .B(n335), .A(n337), .Y(n336) );
  INVX1 U216 ( .A(n349), .Y(n363) );
  AND2XL U217 ( .A(n391), .B(ps_ptr[3]), .Y(N1034) );
  INVXL U218 ( .A(stop), .Y(n302) );
  XNOR3X1 U219 ( .A(N1505), .B(N1503), .C(sub_395_S2_I9_aco_carry[4]), .Y(n396) );
  XNOR3X1 U220 ( .A(N1669), .B(N1667), .C(sub_395_S2_I13_aco_carry[4]), .Y(
        n392) );
  AND2X1 U221 ( .A(n651), .B(n640), .Y(n52) );
  AND2X1 U222 ( .A(n613), .B(n612), .Y(n53) );
  AND2X1 U223 ( .A(n655), .B(n654), .Y(n54) );
  XOR2X1 U224 ( .A(n165), .B(sub_395_S2_I13_aco_carry[2]), .Y(n407) );
  INVX1 U225 ( .A(N1665), .Y(n165) );
  INVX1 U226 ( .A(N1307), .Y(n722) );
  AND2X1 U227 ( .A(n664), .B(n663), .Y(n55) );
  AND2X1 U228 ( .A(n659), .B(n658), .Y(n56) );
  NOR2X1 U229 ( .A(n726), .B(N1305), .Y(n503) );
  INVX1 U230 ( .A(n591), .Y(n680) );
  INVX1 U231 ( .A(n590), .Y(n679) );
  INVX1 U232 ( .A(N1386), .Y(n716) );
  INVX1 U233 ( .A(N1714), .Y(n681) );
  XOR2X1 U234 ( .A(n157), .B(sub_395_S2_I9_aco_carry[2]), .Y(n411) );
  INVX1 U235 ( .A(N1501), .Y(n157) );
  XNOR2XL U236 ( .A(N1666), .B(sub_395_S2_I13_aco_carry[3]), .Y(n401) );
  XOR2X1 U237 ( .A(n417), .B(N1664), .Y(n211) );
  XOR2X1 U238 ( .A(n414), .B(N1500), .Y(n208) );
  NAND21X1 U239 ( .B(n60), .A(n192), .Y(n123) );
  NAND21X1 U240 ( .B(n122), .A(n187), .Y(n133) );
  INVX1 U241 ( .A(N1717), .Y(n677) );
  INVX1 U242 ( .A(N1389), .Y(n712) );
  INVX1 U243 ( .A(n393), .Y(n695) );
  INVX1 U244 ( .A(n406), .Y(n689) );
  INVX1 U245 ( .A(n135), .Y(n673) );
  NAND2X1 U246 ( .A(N1305), .B(n726), .Y(n505) );
  NAND2X1 U247 ( .A(n410), .B(n406), .Y(n578) );
  NAND2X1 U248 ( .A(n410), .B(n689), .Y(n577) );
  NOR2X1 U249 ( .A(n689), .B(n410), .Y(n575) );
  NOR2X1 U250 ( .A(n406), .B(n410), .Y(n576) );
  INVX1 U251 ( .A(n482), .Y(n715) );
  INVX1 U252 ( .A(n506), .Y(n725) );
  INVX1 U253 ( .A(n481), .Y(n714) );
  INVX1 U254 ( .A(N1222), .Y(n736) );
  INVX1 U255 ( .A(N1716), .Y(n678) );
  AO21X1 U256 ( .B(n132), .C(n131), .A(n148), .Y(N1838) );
  AO21X1 U257 ( .B(n123), .C(n122), .A(n121), .Y(N1756) );
  AO21X1 U258 ( .B(n193), .C(n192), .A(n191), .Y(N1837) );
  XNOR2XL U259 ( .A(N1502), .B(sub_395_S2_I9_aco_carry[3]), .Y(n404) );
  XNOR2XL U260 ( .A(N1625), .B(sub_395_S2_I12_aco_carry[3]), .Y(n403) );
  NAND21X1 U261 ( .B(n125), .A(n189), .Y(n138) );
  INVX1 U262 ( .A(N1755), .Y(n676) );
  NAND2X1 U263 ( .A(n409), .B(n405), .Y(n530) );
  NAND2X1 U264 ( .A(N1756), .B(N1755), .Y(n620) );
  NAND2X1 U265 ( .A(n409), .B(n210), .Y(n529) );
  NOR2X1 U266 ( .A(N1222), .B(N1223), .Y(n456) );
  NOR2X1 U267 ( .A(n736), .B(N1223), .Y(n455) );
  INVX1 U268 ( .A(n131), .Y(n191) );
  NOR2X1 U269 ( .A(n210), .B(n409), .Y(n527) );
  NOR2X1 U270 ( .A(n405), .B(n409), .Y(n528) );
  NOR2X1 U271 ( .A(N1755), .B(N1756), .Y(n618) );
  NOR2X1 U272 ( .A(n672), .B(N1797), .Y(n631) );
  NAND21X1 U273 ( .B(n137), .A(n124), .Y(n136) );
  NAND21X1 U274 ( .B(n61), .A(n193), .Y(n665) );
  XNOR2XL U275 ( .A(N1461), .B(sub_395_S2_I8_aco_carry[3]), .Y(n402) );
  INVX1 U276 ( .A(n209), .Y(N1550) );
  NAND2XL U277 ( .A(N1223), .B(N1222), .Y(n458) );
  NAND2X1 U278 ( .A(N1223), .B(n736), .Y(n457) );
  NAND2X1 U279 ( .A(N1797), .B(n672), .Y(n633) );
  INVX1 U280 ( .A(n634), .Y(n671) );
  INVX1 U281 ( .A(n554), .Y(n698) );
  INVX1 U282 ( .A(n553), .Y(n697) );
  AOI21AX1 U283 ( .B(n138), .C(n137), .A(n136), .Y(n57) );
  INVX1 U284 ( .A(n128), .Y(n132) );
  INVX1 U285 ( .A(n147), .Y(n146) );
  INVX1 U286 ( .A(n410), .Y(n161) );
  INVX1 U287 ( .A(n409), .Y(n164) );
  AO21X1 U288 ( .B(N1462), .C(n413), .A(n107), .Y(sub_395_S2_I8_aco_carry[5])
         );
  OA21X1 U289 ( .B(N1462), .C(n413), .A(sub_395_S2_I8_aco_carry[4]), .Y(n107)
         );
  OAI21BBX1 U290 ( .A(N1667), .B(n417), .C(n58), .Y(
        sub_395_S2_I13_aco_carry[5]) );
  OAI21X1 U291 ( .B(N1667), .C(n417), .A(sub_395_S2_I13_aco_carry[4]), .Y(n58)
         );
  AO21X1 U292 ( .B(N1503), .C(n414), .A(n106), .Y(sub_395_S2_I9_aco_carry[5])
         );
  OA21X1 U293 ( .B(N1503), .C(n414), .A(sub_395_S2_I9_aco_carry[4]), .Y(n106)
         );
  AO21X1 U294 ( .B(N1626), .C(n416), .A(n108), .Y(sub_395_S2_I12_aco_carry[5])
         );
  OA21X1 U295 ( .B(N1626), .C(n416), .A(sub_395_S2_I12_aco_carry[4]), .Y(n108)
         );
  AO21XL U296 ( .B(n225), .C(n224), .A(n275), .Y(n227) );
  AOI31XL U297 ( .A(n359), .B(n360), .C(n358), .D(n281), .Y(n228) );
  AOI221XL U298 ( .A(n316), .B(N1345), .C(n312), .D(N1222), .E(n400), .Y(n399)
         );
  AOI22X1 U299 ( .A(n85), .B(n343), .C(n313), .D(N1386), .Y(n398) );
  AOI22XL U300 ( .A(n314), .B(N1263), .C(n315), .D(N1181), .Y(n397) );
  AOI21XL U301 ( .B(n240), .C(n239), .A(n275), .Y(n59) );
  BUFX3 U302 ( .A(n760), .Y(ps_ptr[2]) );
  INVX1 U303 ( .A(N1756), .Y(n186) );
  OA21X1 U304 ( .B(n171), .C(n281), .A(n170), .Y(n185) );
  INVX1 U305 ( .A(N1838), .Y(n183) );
  INVX1 U306 ( .A(N1797), .Y(n181) );
  NOR32XL U307 ( .B(n177), .C(n176), .A(n175), .Y(n182) );
  OAI22X1 U308 ( .A(N1217), .B(n297), .C(n296), .D(n295), .Y(n381) );
  OA222X1 U309 ( .A(N1215), .B(n320), .C(n294), .D(n293), .E(n90), .F(n292), 
        .Y(n296) );
  INVXL U310 ( .A(ps_ptr[2]), .Y(n292) );
  OA21XL U311 ( .B(n276), .C(n275), .A(n274), .Y(n277) );
  AND4X1 U312 ( .A(n273), .B(n369), .C(n370), .D(n272), .Y(n276) );
  INVX3 U313 ( .A(n152), .Y(n178) );
  OAI31XL U314 ( .A(n371), .B(n374), .C(n368), .D(n388), .Y(n270) );
  INVXL U315 ( .A(n275), .Y(n388) );
  NAND32X1 U316 ( .B(n352), .C(n351), .A(n2), .Y(n353) );
  INVX1 U317 ( .A(n357), .Y(n366) );
  INVX1 U318 ( .A(n330), .Y(n345) );
  INVX1 U319 ( .A(n348), .Y(n354) );
  NAND21X1 U320 ( .B(n344), .A(n337), .Y(n349) );
  INVX1 U321 ( .A(n344), .Y(n335) );
  INVX1 U322 ( .A(n328), .Y(n332) );
  INVX1 U323 ( .A(n319), .Y(n364) );
  NAND32X1 U324 ( .B(n335), .C(n327), .A(n332), .Y(n319) );
  INVX1 U325 ( .A(n326), .Y(n329) );
  NAND32X1 U326 ( .B(n328), .C(n327), .A(n335), .Y(n350) );
  INVX1 U327 ( .A(n327), .Y(n331) );
  AND2X1 U328 ( .A(n391), .B(ps_ptr[1]), .Y(N1032) );
  INVX1 U329 ( .A(n203), .Y(n177) );
  OA2222XL U330 ( .A(n210), .B(n273), .C(n209), .D(n370), .E(n208), .F(n269), 
        .G(n689), .H(n369), .Y(n213) );
  INVX1 U331 ( .A(n405), .Y(n210) );
  OA222X1 U332 ( .A(n681), .B(n272), .C(n211), .D(n268), .E(n334), .F(n694), 
        .Y(n212) );
  INVX1 U333 ( .A(n422), .Y(n159) );
  AND3X1 U334 ( .A(n376), .B(n377), .C(n375), .Y(n171) );
  AOI221XL U335 ( .A(n316), .B(N1346), .C(n312), .D(N1223), .E(n378), .Y(n377)
         );
  AOI22X1 U336 ( .A(n91), .B(n343), .C(n313), .D(N1387), .Y(n376) );
  AOI22X1 U337 ( .A(n314), .B(N1264), .C(n315), .D(N1182), .Y(n375) );
  NOR2X1 U338 ( .A(n681), .B(N1715), .Y(n588) );
  NOR2X1 U339 ( .A(N1714), .B(N1715), .Y(n589) );
  INVX1 U340 ( .A(N1304), .Y(n726) );
  XNOR3X1 U341 ( .A(N1628), .B(N1626), .C(sub_395_S2_I12_aco_carry[4]), .Y(
        n395) );
  OA2222XL U342 ( .A(n273), .B(n238), .C(n370), .D(n695), .E(n269), .F(n237), 
        .G(n369), .H(n236), .Y(n240) );
  INVX1 U343 ( .A(n395), .Y(n236) );
  INVX1 U344 ( .A(n394), .Y(n238) );
  OA2222XL U345 ( .A(n702), .B(n273), .C(n696), .D(n370), .E(n699), .F(n269), 
        .G(n686), .H(n369), .Y(n225) );
  OA222X1 U346 ( .A(n678), .B(n272), .C(n683), .D(n268), .E(n334), .F(n691), 
        .Y(n224) );
  OA222X1 U347 ( .A(n334), .B(n690), .C(n268), .D(n682), .E(n677), .F(n272), 
        .Y(n239) );
  INVX1 U348 ( .A(N1628), .Y(n416) );
  NAND2X1 U349 ( .A(N1715), .B(n681), .Y(n590) );
  NAND2XL U350 ( .A(N1715), .B(N1714), .Y(n591) );
  NOR2X1 U351 ( .A(N1386), .B(N1387), .Y(n480) );
  NOR2X1 U352 ( .A(N1304), .B(N1305), .Y(n504) );
  NOR2X1 U353 ( .A(n716), .B(N1387), .Y(n479) );
  INVX1 U354 ( .A(n269), .Y(n374) );
  OAI22X1 U355 ( .A(n705), .B(n711), .C(n726), .D(n342), .Y(n400) );
  AOI22X1 U356 ( .A(n314), .B(N1265), .C(n315), .D(N1183), .Y(n358) );
  AOI221XL U357 ( .A(n316), .B(N1348), .C(n312), .D(N1225), .E(n341), .Y(n340)
         );
  OAI22X1 U358 ( .A(n705), .B(n707), .C(n722), .D(n342), .Y(n341) );
  AOI22X1 U359 ( .A(N1217), .B(n343), .C(n313), .D(N1389), .Y(n339) );
  AOI22X1 U360 ( .A(n314), .B(N1266), .C(n315), .D(N1184), .Y(n338) );
  INVX1 U361 ( .A(n342), .Y(n706) );
  INVX1 U362 ( .A(n334), .Y(n368) );
  XNOR3X1 U363 ( .A(N1546), .B(N1544), .C(sub_395_S2_I10_aco_carry[4]), .Y(
        n393) );
  XNOR3X1 U364 ( .A(N1464), .B(N1462), .C(sub_395_S2_I8_aco_carry[4]), .Y(n394) );
  XOR2X1 U365 ( .A(n416), .B(n83), .Y(n406) );
  XOR2X1 U366 ( .A(N1460), .B(sub_395_S2_I12_aco_carry[2]), .Y(n410) );
  XOR3X1 U367 ( .A(n70), .B(n60), .C(n382), .Y(n135) );
  NAND21X1 U368 ( .B(n69), .A(n121), .Y(n382) );
  INVX1 U369 ( .A(N1464), .Y(n413) );
  INVX1 U370 ( .A(N1546), .Y(n415) );
  NAND2XL U371 ( .A(N1387), .B(N1386), .Y(n482) );
  NAND2XL U372 ( .A(N1305), .B(N1304), .Y(n506) );
  NAND2X1 U373 ( .A(N1387), .B(n716), .Y(n481) );
  AOI21X1 U374 ( .B(n111), .C(n70), .A(N1750), .Y(n60) );
  AOI221XL U375 ( .A(n316), .B(N1347), .C(n312), .D(N1224), .E(n361), .Y(n360)
         );
  OAI22X1 U376 ( .A(n705), .B(n708), .C(n723), .D(n342), .Y(n361) );
  AOI22X1 U377 ( .A(n96), .B(n343), .C(n313), .D(N1388), .Y(n359) );
  AOI22X1 U378 ( .A(n77), .B(n343), .C(n313), .D(n77), .Y(n427) );
  XOR2X1 U379 ( .A(n413), .B(n83), .Y(n405) );
  XOR2X1 U380 ( .A(N1296), .B(sub_395_S2_I8_aco_carry[2]), .Y(n409) );
  AO21X1 U381 ( .B(n126), .C(n125), .A(n124), .Y(N1797) );
  AO21X1 U382 ( .B(n60), .C(n188), .A(n187), .Y(N1755) );
  XOR2X1 U383 ( .A(n129), .B(n95), .Y(n147) );
  NAND21X1 U384 ( .B(n127), .A(cs_ptr[2]), .Y(n129) );
  AOI21BX1 U385 ( .C(n129), .B(n96), .A(N1217), .Y(n61) );
  NAND21X1 U386 ( .B(n192), .A(n144), .Y(n131) );
  INVX1 U387 ( .A(N1225), .Y(n732) );
  INVX1 U388 ( .A(N1796), .Y(n672) );
  INVX1 U389 ( .A(n126), .Y(n189) );
  NOR2X1 U390 ( .A(n209), .B(n408), .Y(n551) );
  INVX1 U391 ( .A(n268), .Y(n371) );
  INVX1 U392 ( .A(n144), .Y(n193) );
  INVX1 U393 ( .A(n119), .Y(n190) );
  NAND21X1 U394 ( .B(n120), .A(n136), .Y(n669) );
  XOR2X1 U395 ( .A(n116), .B(n190), .Y(n120) );
  INVX1 U396 ( .A(n114), .Y(n116) );
  XOR2X1 U397 ( .A(n127), .B(n89), .Y(n128) );
  XOR2X1 U398 ( .A(n415), .B(n83), .Y(n209) );
  INVX1 U399 ( .A(n188), .Y(n192) );
  NAND2X1 U400 ( .A(N1797), .B(N1796), .Y(n634) );
  NAND2X1 U401 ( .A(n408), .B(n209), .Y(n553) );
  NAND2X1 U402 ( .A(n408), .B(N1550), .Y(n554) );
  INVX1 U403 ( .A(n112), .Y(n122) );
  AOI21AX1 U404 ( .B(n133), .C(n69), .A(n382), .Y(n62) );
  NOR2X1 U405 ( .A(N1796), .B(N1797), .Y(n632) );
  NOR2X1 U406 ( .A(N1550), .B(n408), .Y(n552) );
  INVX1 U407 ( .A(N1715), .Y(n168) );
  ENOX1 U408 ( .A(n63), .B(n370), .C(N1677), .D(n371), .Y(n372) );
  XOR2X1 U409 ( .A(N1545), .B(sub_395_S2_I10_aco_carry[5]), .Y(n63) );
  INVX1 U410 ( .A(n117), .Y(n137) );
  INVX1 U411 ( .A(n118), .Y(n125) );
  INVX1 U412 ( .A(n369), .Y(n373) );
  INVX1 U413 ( .A(n408), .Y(n163) );
  OAI21BBX1 U414 ( .A(N1544), .B(n415), .C(n64), .Y(
        sub_395_S2_I10_aco_carry[5]) );
  OAI21X1 U415 ( .B(N1544), .C(n415), .A(sub_395_S2_I10_aco_carry[4]), .Y(n64)
         );
  AOI21XL U416 ( .B(n213), .C(n212), .A(n275), .Y(n65) );
  INVX1 U417 ( .A(n155), .Y(n154) );
  NAND32XL U418 ( .B(wr_dacv[13]), .C(n244), .A(n26), .Y(n196) );
  OAI22XL U419 ( .A(ps_ptr[1]), .B(n87), .C(ps_ptr[2]), .D(n93), .Y(n293) );
  INVX1 U420 ( .A(n194), .Y(n254) );
  NAND5XL U421 ( .A(n173), .B(n249), .C(n248), .D(n41), .E(n29), .Y(n231) );
  INVX1 U422 ( .A(n196), .Y(n173) );
  NAND32X1 U423 ( .B(n307), .C(n275), .A(n156), .Y(n281) );
  INVX1 U424 ( .A(n305), .Y(n156) );
  NAND2XL U425 ( .A(n172), .B(n178), .Y(n271) );
  AOI22BXL U426 ( .B(N1795), .A(ps_ptr[0]), .D(n84), .C(ps_ptr[1]), .Y(n294)
         );
  NAND32XL U427 ( .B(wr_dacv[16]), .C(n246), .A(n5), .Y(n247) );
  AOI21BBXL U428 ( .B(n79), .C(ps_ptr[0]), .A(n381), .Y(n298) );
  NAND32XL U429 ( .B(stop), .C(n105), .A(n390), .Y(n660) );
  MUX2X1 U430 ( .D0(busy), .D1(n389), .S(n391), .Y(n390) );
  AOI222XL U431 ( .A(n388), .B(n387), .C(n386), .D(busy), .E(n385), .F(n384), 
        .Y(n389) );
  AND3X1 U432 ( .A(n382), .B(n70), .C(N1750), .Y(n385) );
  NAND32X1 U433 ( .B(n331), .C(n105), .A(n318), .Y(N1002) );
  OA22X1 U434 ( .A(n317), .B(n303), .C(ps_sample), .D(n302), .Y(n318) );
  AND4X1 U435 ( .A(ps_sample), .B(n300), .C(n299), .D(n298), .Y(n317) );
  NAND6XL U436 ( .A(n73), .B(n205), .C(n207), .D(n266), .E(n32), .F(n35), .Y(
        n218) );
  AND3X1 U437 ( .A(n266), .B(n35), .C(n265), .Y(n267) );
  AND3X1 U438 ( .A(n223), .B(n234), .C(n222), .Y(n229) );
  INVX1 U439 ( .A(n174), .Y(n235) );
  NAND43X1 U440 ( .B(n194), .C(n253), .D(n243), .A(n195), .Y(n174) );
  INVX1 U441 ( .A(n255), .Y(n195) );
  OAI211X1 U442 ( .C(n197), .D(n196), .A(n254), .B(n195), .Y(n198) );
  INVX1 U443 ( .A(n347), .Y(n352) );
  AND3X1 U444 ( .A(n367), .B(n366), .C(n365), .Y(N1003) );
  AND2X1 U445 ( .A(n364), .B(n355), .Y(N1012) );
  AND2X1 U446 ( .A(n367), .B(n355), .Y(N1011) );
  OAI32X1 U447 ( .A(n357), .B(n350), .C(n365), .D(n349), .E(n348), .Y(N1013)
         );
  MUX2XL U448 ( .D0(N1215), .D1(ps_ptr[3]), .S(ps_sample), .Y(n351) );
  MUX2XL U449 ( .D0(n85), .D1(ps_ptr[1]), .S(ps_sample), .Y(n328) );
  NAND21X1 U450 ( .B(n105), .A(n291), .Y(n327) );
  MUX2X1 U451 ( .D0(n290), .D1(n283), .S(ps_sample), .Y(n291) );
  AND3X1 U452 ( .A(sampl_begn), .B(n302), .C(n303), .Y(n290) );
  NAND21X1 U453 ( .B(n262), .A(n261), .Y(n203) );
  INVX1 U454 ( .A(n201), .Y(n259) );
  INVX1 U455 ( .A(n219), .Y(n261) );
  INVX1 U456 ( .A(n202), .Y(n217) );
  NAND21X1 U457 ( .B(n260), .A(n259), .Y(n202) );
  INVX1 U458 ( .A(n258), .Y(n205) );
  INVX1 U459 ( .A(n260), .Y(n176) );
  INVX1 U460 ( .A(n262), .Y(n234) );
  NAND2X1 U461 ( .A(sampl_done), .B(srstz), .Y(n322) );
  NOR2X1 U462 ( .A(n322), .B(n759), .Y(N971) );
  NOR2X1 U463 ( .A(n48), .B(n758), .Y(N970) );
  NOR2X1 U464 ( .A(n322), .B(n757), .Y(N969) );
  NOR2X1 U465 ( .A(n48), .B(n756), .Y(N968) );
  NOR2X1 U466 ( .A(n322), .B(n755), .Y(N967) );
  NOR2X1 U467 ( .A(n48), .B(n754), .Y(N966) );
  NOR2X1 U468 ( .A(n322), .B(n753), .Y(N963) );
  NOR2X1 U469 ( .A(n48), .B(n752), .Y(N962) );
  NOR2X1 U470 ( .A(n322), .B(n751), .Y(N961) );
  NOR2X1 U471 ( .A(n48), .B(n750), .Y(N960) );
  NOR2X1 U472 ( .A(n322), .B(n749), .Y(N959) );
  NOR2X1 U473 ( .A(n48), .B(n748), .Y(N958) );
  NOR2X1 U474 ( .A(n322), .B(n747), .Y(N957) );
  NOR2X1 U475 ( .A(n48), .B(n746), .Y(N956) );
  NOR32XL U476 ( .B(n421), .C(n419), .A(n420), .Y(n422) );
  NAND31X1 U477 ( .C(n431), .A(n432), .B(n430), .Y(n434) );
  NAND21X1 U478 ( .B(n159), .A(n424), .Y(n370) );
  NOR21XL U479 ( .B(n437), .A(n438), .Y(n343) );
  NAND32X1 U480 ( .B(n160), .C(n159), .A(n158), .Y(n269) );
  INVX1 U481 ( .A(n424), .Y(n158) );
  INVX1 U482 ( .A(n423), .Y(n160) );
  NAND32X1 U483 ( .B(n423), .C(n424), .A(n422), .Y(n305) );
  NAND21X1 U484 ( .B(n305), .A(n307), .Y(n273) );
  AND2X1 U485 ( .A(n425), .B(n418), .Y(n66) );
  AND2X1 U486 ( .A(n437), .B(n438), .Y(n315) );
  NAND3X1 U487 ( .A(n419), .B(n420), .C(n421), .Y(n334) );
  INVX1 U488 ( .A(n98), .Y(cs_ptr[3]) );
  INVX1 U489 ( .A(n92), .Y(cs_ptr[2]) );
  INVX1 U490 ( .A(n104), .Y(cs_ptr[4]) );
  INVX1 U491 ( .A(n99), .Y(n95) );
  INVX1 U492 ( .A(n87), .Y(n83) );
  INVX1 U493 ( .A(n92), .Y(n89) );
  INVX1 U494 ( .A(n80), .Y(n76) );
  NOR2X1 U495 ( .A(n301), .B(n583), .Y(n421) );
  INVX1 U496 ( .A(n92), .Y(n90) );
  NOR2X1 U497 ( .A(n311), .B(n436), .Y(n432) );
  INVX1 U498 ( .A(n79), .Y(n77) );
  INVX1 U499 ( .A(n87), .Y(n85) );
  INVX1 U500 ( .A(n93), .Y(n91) );
  NOR3XL U501 ( .A(n434), .B(n435), .C(n433), .Y(n437) );
  INVX1 U502 ( .A(n79), .Y(n78) );
  AND2X1 U503 ( .A(n657), .B(n656), .Y(n67) );
  AND2X1 U504 ( .A(n653), .B(n652), .Y(n68) );
  NOR21XL U505 ( .B(n432), .A(n430), .Y(n316) );
  NOR21XL U506 ( .B(n435), .A(n434), .Y(n314) );
  NAND21X1 U507 ( .B(n419), .A(n421), .Y(n369) );
  NAND21X1 U508 ( .B(n301), .A(n583), .Y(n268) );
  AO22X1 U509 ( .A(n311), .B(N1428), .C(N1305), .D(n706), .Y(n378) );
  NOR31X1 U510 ( .C(n433), .A(n434), .B(n435), .Y(n312) );
  NAND3X1 U511 ( .A(n430), .B(n431), .C(n432), .Y(n342) );
  INVX1 U512 ( .A(n104), .Y(n101) );
  INVX1 U513 ( .A(n104), .Y(n102) );
  INVX1 U514 ( .A(n86), .Y(n84) );
  INVX1 U515 ( .A(n99), .Y(n96) );
  INVX1 U516 ( .A(n311), .Y(n705) );
  INVX1 U517 ( .A(n301), .Y(n272) );
  INVX1 U518 ( .A(n98), .Y(n97) );
  XNOR2XL U519 ( .A(n98), .B(add_394_I15_carry_3_), .Y(n69) );
  AND2X1 U520 ( .A(n436), .B(n705), .Y(n313) );
  INVX1 U521 ( .A(n87), .Y(cs_ptr[1]) );
  INVX1 U522 ( .A(n80), .Y(cs_ptr[0]) );
  XNOR2XL U523 ( .A(n103), .B(add_394_I15_carry_4_), .Y(n70) );
  AND2X1 U524 ( .A(n662), .B(n661), .Y(n71) );
  XOR2X1 U525 ( .A(n92), .B(sub_395_S2_I10_aco_carry[2]), .Y(n408) );
  AO21X1 U526 ( .B(n190), .C(n87), .A(n189), .Y(N1796) );
  XOR2X1 U527 ( .A(n92), .B(add_394_I15_carry_2_), .Y(n112) );
  OAI21BBX1 U528 ( .A(n86), .B(n81), .C(n127), .Y(n188) );
  NAND21X1 U529 ( .B(n79), .A(cs_ptr[1]), .Y(n127) );
  XOR2X1 U530 ( .A(n103), .B(add_394_I16_carry[4]), .Y(n114) );
  NAND21X1 U531 ( .B(n87), .A(n119), .Y(n126) );
  OAI22X1 U532 ( .A(n103), .B(n115), .C(n114), .D(n113), .Y(n119) );
  INVX1 U533 ( .A(add_394_I16_carry[4]), .Y(n115) );
  AND3X1 U534 ( .A(n117), .B(n83), .C(n118), .Y(n113) );
  OAI22X1 U535 ( .A(n103), .B(n98), .C(n130), .D(n61), .Y(n144) );
  AND3X1 U536 ( .A(n128), .B(n188), .C(n147), .Y(n130) );
  AOI221XL U537 ( .A(n316), .B(n80), .C(n312), .D(n77), .E(n429), .Y(n428) );
  OAI22X1 U538 ( .A(n705), .B(n77), .C(n81), .D(n342), .Y(n429) );
  XOR2X1 U539 ( .A(n98), .B(add_394_I16_carry[3]), .Y(n117) );
  XOR2X1 U540 ( .A(n86), .B(cs_ptr[2]), .Y(n118) );
  XOR2X1 U541 ( .A(n98), .B(sub_395_S2_I10_aco_carry[3]), .Y(n696) );
  OAI211X1 U542 ( .C(n304), .D(n305), .A(n380), .B(n379), .Y(n387) );
  AOI22X1 U543 ( .A(N1595), .B(n368), .C(N1718), .D(n301), .Y(n380) );
  AOI221XL U544 ( .A(N1513), .B(n374), .C(N1636), .D(n373), .E(n372), .Y(n379)
         );
  AOI22X1 U545 ( .A(n412), .B(n306), .C(N1472), .D(n307), .Y(n304) );
  NAND3X1 U546 ( .A(n308), .B(n309), .C(n310), .Y(n306) );
  AOI22X1 U547 ( .A(N1390), .B(n313), .C(N1267), .D(n314), .Y(n309) );
  AOI222XL U548 ( .A(N1431), .B(n311), .C(N1226), .D(n312), .E(N1308), .F(n706), .Y(n310) );
  AOI22X1 U549 ( .A(N1185), .B(n315), .C(N1349), .D(n316), .Y(n308) );
  INVX1 U550 ( .A(n307), .Y(n412) );
  MUX2IX1 U551 ( .D0(n245), .D1(n5), .S(cs_ptr[0]), .Y(n72) );
  INVX1 U552 ( .A(sampl_done), .Y(n303) );
  AND2X1 U553 ( .A(n98), .B(n103), .Y(n323) );
  NAND4X1 U554 ( .A(n746), .B(n754), .C(n755), .D(n756), .Y(n287) );
  NOR4XL U555 ( .A(n284), .B(n285), .C(n286), .D(n287), .Y(sh_hold) );
  NAND4X1 U556 ( .A(n747), .B(n748), .C(n749), .D(n750), .Y(n285) );
  NAND4X1 U557 ( .A(n751), .B(n752), .C(n289), .D(n753), .Y(n284) );
  OR2XL U558 ( .A(wr_dacv[10]), .B(n19), .Y(n194) );
  OR2XL U559 ( .A(wr_dacv[12]), .B(n25), .Y(n244) );
  OAI211X1 U560 ( .C(n282), .D(n281), .A(n280), .B(n279), .Y(ps_ptr[0]) );
  AND3X1 U561 ( .A(n427), .B(n428), .C(n426), .Y(n282) );
  OAI31XL U562 ( .A(n267), .B(n33), .C(wr_dacv[1]), .D(n73), .Y(n280) );
  MUX2X1 U563 ( .D0(n278), .D1(n277), .S(cs_ptr[0]), .Y(n279) );
  NAND43X1 U564 ( .B(wr_dacv[16]), .C(wr_dacv[17]), .D(n7), .A(n245), .Y(n221)
         );
  OR2XL U565 ( .A(wr_dacv[9]), .B(n16), .Y(n253) );
  OR2XL U566 ( .A(wr_dacv[11]), .B(n22), .Y(n255) );
  AND4X1 U567 ( .A(n200), .B(n199), .C(n198), .D(n38), .Y(n204) );
  OAI21AX1 U568 ( .B(r_loop), .C(n381), .A(r_semi), .Y(n386) );
  OAI211X1 U569 ( .C(n252), .D(n251), .A(n250), .B(n26), .Y(n256) );
  INVXL U570 ( .A(wr_dacv[13]), .Y(n250) );
  NAND21X1 U571 ( .B(n42), .A(n249), .Y(n251) );
  AND3X1 U572 ( .A(n248), .B(n29), .C(n247), .Y(n252) );
  NAND21X1 U573 ( .B(n40), .A(n199), .Y(n243) );
  AO21X1 U574 ( .B(ps_md4ch), .C(n325), .A(n324), .Y(n347) );
  MUX2XL U575 ( .D0(n90), .D1(ps_ptr[2]), .S(ps_sample), .Y(n324) );
  MUX2BXL U576 ( .D0(n323), .D1(n321), .S(ps_sample), .Y(n325) );
  AO21X1 U577 ( .B(r_comp_swtch), .C(n356), .A(n354), .Y(n355) );
  OR2X1 U578 ( .A(wr_dacv[7]), .B(r_dac_en[7]), .Y(n262) );
  OR2X1 U579 ( .A(wr_dacv[5]), .B(r_dac_en[5]), .Y(n260) );
  OR2X1 U580 ( .A(wr_dacv[6]), .B(r_dac_en[6]), .Y(n219) );
  OR2X1 U581 ( .A(wr_dacv[4]), .B(r_dac_en[4]), .Y(n201) );
  OR2X1 U582 ( .A(wr_dacv[3]), .B(n13), .Y(n258) );
  NOR21XL U583 ( .B(pos_dacis[17]), .A(n322), .Y(N973) );
  NOR21XL U584 ( .B(pos_dacis[16]), .A(n48), .Y(N972) );
  NOR21XL U585 ( .B(pos_dacis[8]), .A(n322), .Y(N964) );
  NOR21XL U586 ( .B(pos_dacis[9]), .A(n48), .Y(N965) );
  INVX1 U587 ( .A(cs_mux_5_), .Y(busy) );
  OR2X1 U588 ( .A(neg_dacis[11]), .B(pos_dacis[11]), .Y(app_dacis[11]) );
  OR2X1 U589 ( .A(neg_dacis[6]), .B(pos_dacis[6]), .Y(app_dacis[6]) );
  OR2X1 U590 ( .A(neg_dacis[7]), .B(pos_dacis[7]), .Y(app_dacis[7]) );
  OR2X1 U591 ( .A(neg_dacis[16]), .B(pos_dacis[16]), .Y(app_dacis[16]) );
  OR2X1 U592 ( .A(neg_dacis[0]), .B(pos_dacis[0]), .Y(app_dacis[0]) );
  OR2X1 U593 ( .A(neg_dacis[14]), .B(pos_dacis[14]), .Y(app_dacis[14]) );
  OR2X1 U594 ( .A(neg_dacis[12]), .B(pos_dacis[12]), .Y(app_dacis[12]) );
  OR2X1 U595 ( .A(neg_dacis[15]), .B(pos_dacis[15]), .Y(app_dacis[15]) );
  OR2X1 U596 ( .A(neg_dacis[5]), .B(pos_dacis[5]), .Y(app_dacis[5]) );
  OR2X1 U597 ( .A(neg_dacis[17]), .B(pos_dacis[17]), .Y(app_dacis[17]) );
  OR2X1 U598 ( .A(neg_dacis[2]), .B(pos_dacis[2]), .Y(app_dacis[2]) );
  OR2X1 U599 ( .A(neg_dacis[3]), .B(pos_dacis[3]), .Y(app_dacis[3]) );
  OR2X1 U600 ( .A(neg_dacis[13]), .B(pos_dacis[13]), .Y(app_dacis[13]) );
  OR2X1 U601 ( .A(neg_dacis[10]), .B(pos_dacis[10]), .Y(app_dacis[10]) );
  OR2X1 U602 ( .A(neg_dacis[8]), .B(pos_dacis[8]), .Y(app_dacis[8]) );
  OR2X1 U603 ( .A(neg_dacis[4]), .B(pos_dacis[4]), .Y(app_dacis[4]) );
  OR2X1 U604 ( .A(neg_dacis[1]), .B(pos_dacis[1]), .Y(app_dacis[1]) );
  OR2X1 U605 ( .A(neg_dacis[9]), .B(pos_dacis[9]), .Y(app_dacis[9]) );
  INVX1 U606 ( .A(pos_dacis[14]), .Y(n758) );
  INVX1 U607 ( .A(pos_dacis[12]), .Y(n756) );
  INVX1 U608 ( .A(pos_dacis[15]), .Y(n759) );
  INVX1 U609 ( .A(pos_dacis[6]), .Y(n752) );
  INVX1 U610 ( .A(pos_dacis[7]), .Y(n753) );
  INVX1 U611 ( .A(pos_dacis[5]), .Y(n751) );
  INVX1 U612 ( .A(pos_dacis[4]), .Y(n750) );
  INVX1 U613 ( .A(pos_dacis[3]), .Y(n749) );
  INVX1 U614 ( .A(pos_dacis[10]), .Y(n754) );
  INVX1 U615 ( .A(pos_dacis[2]), .Y(n748) );
  INVX1 U616 ( .A(pos_dacis[0]), .Y(n746) );
  INVX1 U617 ( .A(pos_dacis[13]), .Y(n757) );
  INVX1 U618 ( .A(pos_dacis[11]), .Y(n755) );
  INVX1 U619 ( .A(pos_dacis[1]), .Y(n747) );
  OAI22X1 U620 ( .A(n487), .B(n77), .C(n81), .D(n488), .Y(n311) );
  AOI222XL U621 ( .A(N1430), .B(r_dac_en[17]), .C(n496), .D(n708), .E(N1429), 
        .F(n497), .Y(n487) );
  AOI222XL U622 ( .A(N1430), .B(n6), .C(n489), .D(n708), .E(N1429), .F(n490), 
        .Y(n488) );
  AO2222XL U623 ( .A(n710), .B(n30), .C(n709), .D(n27), .E(n491), .F(n21), .G(
        n492), .H(n15), .Y(n497) );
  OAI22X1 U624 ( .A(n584), .B(n79), .C(n78), .D(n585), .Y(n301) );
  AOI222XL U625 ( .A(N1717), .B(r_dac_en[17]), .C(n593), .D(n678), .E(N1716), 
        .F(n594), .Y(n584) );
  AOI222XL U626 ( .A(N1717), .B(n6), .C(n586), .D(n678), .E(N1716), .F(n587), 
        .Y(n585) );
  AO2222XL U627 ( .A(n680), .B(n30), .C(n679), .D(n27), .E(n588), .F(n21), .G(
        n589), .H(n15), .Y(n594) );
  AO2222XL U628 ( .A(n693), .B(n43), .C(n692), .D(n25), .E(n563), .F(n19), .G(
        n564), .H(n40), .Y(n562) );
  OAI22AX1 U629 ( .D(n79), .C(n535), .A(n80), .B(n536), .Y(n423) );
  AOI222XL U630 ( .A(n396), .B(n4), .C(n544), .D(n699), .E(n404), .F(n545), 
        .Y(n535) );
  AOI222XL U631 ( .A(n396), .B(n7), .C(n537), .D(n699), .E(n404), .F(n538), 
        .Y(n536) );
  AO2222XL U632 ( .A(n701), .B(n31), .C(n700), .D(n28), .E(n539), .F(n22), .G(
        n540), .H(n16), .Y(n545) );
  OAI22AX1 U633 ( .D(n81), .C(n596), .A(n81), .B(n597), .Y(n583) );
  AOI222XL U634 ( .A(n392), .B(r_dac_en[17]), .C(n605), .D(n683), .E(n401), 
        .F(n606), .Y(n596) );
  AOI222XL U635 ( .A(n392), .B(n7), .C(n598), .D(n683), .E(n401), .F(n599), 
        .Y(n597) );
  AO2222XL U636 ( .A(n685), .B(n31), .C(n684), .D(n28), .E(n600), .F(n22), .G(
        n601), .H(n16), .Y(n606) );
  OAI22X1 U637 ( .A(n559), .B(n77), .C(n81), .D(n560), .Y(n420) );
  AOI222XL U638 ( .A(N1594), .B(n4), .C(n568), .D(n691), .E(N1593), .F(n569), 
        .Y(n559) );
  AOI222XL U639 ( .A(N1594), .B(n7), .C(n561), .D(n691), .E(N1593), .F(n562), 
        .Y(n560) );
  AO2222XL U640 ( .A(n693), .B(n30), .C(n692), .D(n27), .E(n563), .F(n21), .G(
        n564), .H(n15), .Y(n569) );
  OAI221X1 U641 ( .A(n45), .B(n541), .C(n47), .D(n542), .E(n543), .Y(n537) );
  AOI32X1 U642 ( .A(n10), .B(n237), .C(n540), .D(n539), .E(n37), .Y(n543) );
  OAI221X1 U643 ( .A(n44), .B(n541), .C(n46), .D(n542), .E(n546), .Y(n544) );
  AOI32X1 U644 ( .A(n34), .B(n237), .C(n540), .D(n539), .E(n13), .Y(n546) );
  OAI221X1 U645 ( .A(n745), .B(n602), .C(n743), .D(n603), .E(n604), .Y(n598)
         );
  AOI32X1 U646 ( .A(n10), .B(n682), .C(n601), .D(n600), .E(n37), .Y(n604) );
  OAI221X1 U647 ( .A(n745), .B(n565), .C(n743), .D(n566), .E(n567), .Y(n561)
         );
  AOI32X1 U648 ( .A(n10), .B(n690), .C(n564), .D(n563), .E(n37), .Y(n567) );
  OAI221X1 U649 ( .A(n745), .B(n493), .C(n743), .D(n494), .E(n495), .Y(n489)
         );
  AOI32X1 U650 ( .A(n9), .B(n707), .C(n492), .D(n491), .E(n36), .Y(n495) );
  OAI221X1 U651 ( .A(n744), .B(n493), .C(n742), .D(n494), .E(n498), .Y(n496)
         );
  AOI32X1 U652 ( .A(n33), .B(n707), .C(n492), .D(n491), .E(n12), .Y(n498) );
  OAI221X1 U653 ( .A(n745), .B(n590), .C(n743), .D(n591), .E(n592), .Y(n586)
         );
  AOI32X1 U654 ( .A(n9), .B(n677), .C(n589), .D(n588), .E(n36), .Y(n592) );
  OAI221X1 U655 ( .A(n744), .B(n590), .C(n742), .D(n591), .E(n595), .Y(n593)
         );
  AOI32X1 U656 ( .A(n33), .B(n677), .C(n589), .D(n588), .E(n12), .Y(n595) );
  OAI221X1 U657 ( .A(n744), .B(n565), .C(n742), .D(n566), .E(n570), .Y(n568)
         );
  AOI32X1 U658 ( .A(n33), .B(n690), .C(n564), .D(n563), .E(n12), .Y(n570) );
  OAI221X1 U659 ( .A(n744), .B(n602), .C(n742), .D(n603), .E(n607), .Y(n605)
         );
  AOI32X1 U660 ( .A(n34), .B(n682), .C(n601), .D(n600), .E(n13), .Y(n607) );
  INVX1 U661 ( .A(N1705), .Y(n87) );
  INVX1 U662 ( .A(N1217), .Y(n104) );
  INVX1 U663 ( .A(N1215), .Y(n98) );
  INVX1 U664 ( .A(N1542), .Y(n93) );
  INVX1 U665 ( .A(N1215), .Y(n99) );
  INVX1 U666 ( .A(N1542), .Y(n92) );
  INVX1 U667 ( .A(N1795), .Y(n79) );
  INVX1 U668 ( .A(N1795), .Y(n80) );
  AO2222XL U669 ( .A(n720), .B(n42), .C(n719), .D(n24), .E(n467), .F(n18), .G(
        n468), .H(n39), .Y(n466) );
  AO2222XL U670 ( .A(n710), .B(n42), .C(n709), .D(n24), .E(n491), .F(n18), .G(
        n492), .H(n39), .Y(n490) );
  AO2222XL U671 ( .A(n680), .B(n42), .C(n679), .D(n24), .E(n588), .F(n18), .G(
        n589), .H(n39), .Y(n587) );
  AO2222XL U672 ( .A(n720), .B(n31), .C(n719), .D(n28), .E(n467), .F(n22), .G(
        n468), .H(n16), .Y(n473) );
  EORX1 U673 ( .A(n463), .B(n79), .C(n79), .D(n464), .Y(n430) );
  AOI222XL U674 ( .A(N1348), .B(n6), .C(n465), .D(n718), .E(N1347), .F(n466), 
        .Y(n464) );
  AO222X1 U675 ( .A(N1348), .B(n4), .C(n472), .D(n718), .E(N1347), .F(n473), 
        .Y(n463) );
  INVX1 U676 ( .A(N1347), .Y(n718) );
  OAI22AX1 U677 ( .D(n81), .C(n439), .A(n81), .B(n440), .Y(n438) );
  AOI222XL U678 ( .A(N1184), .B(n4), .C(n448), .D(n738), .E(N1183), .F(n449), 
        .Y(n439) );
  AOI222XL U679 ( .A(N1184), .B(n6), .C(n441), .D(n738), .E(N1183), .F(n442), 
        .Y(n440) );
  INVX1 U680 ( .A(N1183), .Y(n738) );
  OAI22AX1 U681 ( .D(n78), .C(n475), .A(n78), .B(n476), .Y(n436) );
  AOI222XL U682 ( .A(N1389), .B(r_dac_en[17]), .C(n484), .D(n713), .E(N1388), 
        .F(n485), .Y(n475) );
  AOI222XL U683 ( .A(N1389), .B(n7), .C(n477), .D(n713), .E(N1388), .F(n478), 
        .Y(n476) );
  INVX1 U684 ( .A(N1388), .Y(n713) );
  OAI22AX1 U685 ( .D(n81), .C(n511), .A(n81), .B(n512), .Y(n435) );
  AOI222XL U686 ( .A(N1266), .B(n4), .C(n520), .D(n728), .E(N1265), .F(n521), 
        .Y(n511) );
  AOI222XL U687 ( .A(N1266), .B(n6), .C(n513), .D(n728), .E(N1265), .F(n514), 
        .Y(n512) );
  INVX1 U688 ( .A(N1265), .Y(n728) );
  EORX1 U689 ( .A(n571), .B(n76), .C(n77), .D(n572), .Y(n419) );
  AOI222XL U690 ( .A(n395), .B(n6), .C(n573), .D(n686), .E(n403), .F(n574), 
        .Y(n572) );
  AO222X1 U691 ( .A(n395), .B(n4), .C(n580), .D(n686), .E(n403), .F(n581), .Y(
        n571) );
  AO2222XL U692 ( .A(n688), .B(n43), .C(n687), .D(n25), .E(n575), .F(n19), .G(
        n576), .H(n40), .Y(n574) );
  OAI22X1 U693 ( .A(n499), .B(n79), .C(n78), .D(n500), .Y(n431) );
  AOI222XL U694 ( .A(N1307), .B(r_dac_en[17]), .C(n508), .D(n723), .E(N1306), 
        .F(n509), .Y(n499) );
  AOI222XL U695 ( .A(N1307), .B(n7), .C(n501), .D(n723), .E(N1306), .F(n502), 
        .Y(n500) );
  AO2222XL U696 ( .A(n725), .B(n30), .C(n724), .D(n27), .E(n503), .F(n21), .G(
        n504), .H(n15), .Y(n509) );
  OAI221X1 U697 ( .A(n745), .B(n577), .C(n743), .D(n578), .E(n579), .Y(n573)
         );
  AOI32X1 U698 ( .A(n9), .B(n236), .C(n576), .D(n575), .E(n36), .Y(n579) );
  OAI221X1 U699 ( .A(n45), .B(n445), .C(n47), .D(n446), .E(n447), .Y(n441) );
  AOI32X1 U700 ( .A(n9), .B(n737), .C(n444), .D(n443), .E(n36), .Y(n447) );
  OAI221X1 U701 ( .A(n745), .B(n505), .C(n743), .D(n506), .E(n507), .Y(n501)
         );
  AOI32X1 U702 ( .A(n10), .B(n722), .C(n504), .D(n503), .E(n37), .Y(n507) );
  OAI221X1 U703 ( .A(n744), .B(n505), .C(n742), .D(n506), .E(n510), .Y(n508)
         );
  AOI32X1 U704 ( .A(n33), .B(n722), .C(n504), .D(n503), .E(n12), .Y(n510) );
  OAI221X1 U705 ( .A(n745), .B(n481), .C(n743), .D(n482), .E(n483), .Y(n477)
         );
  AOI32X1 U706 ( .A(n10), .B(n712), .C(n480), .D(n479), .E(n37), .Y(n483) );
  OAI221X1 U707 ( .A(n745), .B(n469), .C(n743), .D(n470), .E(n471), .Y(n465)
         );
  AOI32X1 U708 ( .A(n9), .B(n717), .C(n468), .D(n467), .E(n36), .Y(n471) );
  OAI221X1 U709 ( .A(n745), .B(n517), .C(n743), .D(n518), .E(n519), .Y(n513)
         );
  AOI32X1 U710 ( .A(n9), .B(n727), .C(n516), .D(n515), .E(n36), .Y(n519) );
  OAI221X1 U711 ( .A(n744), .B(n577), .C(n742), .D(n578), .E(n582), .Y(n580)
         );
  AOI32X1 U712 ( .A(n34), .B(n236), .C(n576), .D(n575), .E(n13), .Y(n582) );
  OAI221X1 U713 ( .A(n744), .B(n469), .C(n742), .D(n470), .E(n474), .Y(n472)
         );
  AOI32X1 U714 ( .A(n34), .B(n717), .C(n468), .D(n467), .E(n13), .Y(n474) );
  OAI221X1 U715 ( .A(n44), .B(n445), .C(n46), .D(n446), .E(n450), .Y(n448) );
  AOI32X1 U716 ( .A(n33), .B(n737), .C(n444), .D(n443), .E(n12), .Y(n450) );
  OAI221X1 U717 ( .A(n744), .B(n481), .C(n742), .D(n482), .E(n486), .Y(n484)
         );
  AOI32X1 U718 ( .A(n34), .B(n712), .C(n480), .D(n479), .E(n13), .Y(n486) );
  OAI221X1 U719 ( .A(n744), .B(n517), .C(n742), .D(n518), .E(n522), .Y(n520)
         );
  AOI32X1 U720 ( .A(n33), .B(n727), .C(n516), .D(n515), .E(n12), .Y(n522) );
  INVX1 U721 ( .A(N1705), .Y(n86) );
  OAI22AX1 U722 ( .D(n78), .C(n523), .A(N1795), .B(n524), .Y(n307) );
  AOI222XL U723 ( .A(n394), .B(n4), .C(n532), .D(n702), .E(n402), .F(n533), 
        .Y(n523) );
  AOI222XL U724 ( .A(n394), .B(n7), .C(n525), .D(n702), .E(n402), .F(n526), 
        .Y(n524) );
  AO2222XL U725 ( .A(n704), .B(n31), .C(n703), .D(n28), .E(n527), .F(n22), .G(
        n528), .H(n16), .Y(n533) );
  AO21X1 U726 ( .B(n135), .C(n72), .A(n134), .Y(n155) );
  MUX4X1 U727 ( .D0(n623), .D1(n622), .D2(n616), .D3(n615), .S0(n62), .S1(
        cs_ptr[0]), .Y(n134) );
  AO2222XL U728 ( .A(n675), .B(n43), .C(n674), .D(n25), .E(n617), .F(n19), .G(
        n618), .H(n40), .Y(n616) );
  AO2222XL U729 ( .A(n675), .B(n31), .C(n674), .D(n28), .E(n617), .F(n22), .G(
        n618), .H(n16), .Y(n623) );
  OAI22AX1 U730 ( .D(n78), .C(n547), .A(n78), .B(n548), .Y(n424) );
  AOI222XL U731 ( .A(n393), .B(n4), .C(n556), .D(n696), .E(N1552), .F(n557), 
        .Y(n547) );
  AOI222XL U732 ( .A(n393), .B(n6), .C(n549), .D(n696), .E(N1552), .F(n550), 
        .Y(n548) );
  INVX1 U733 ( .A(n696), .Y(N1552) );
  AO2222XL U734 ( .A(n701), .B(n43), .C(n700), .D(n25), .E(n539), .F(n19), .G(
        n540), .H(n40), .Y(n538) );
  AO2222XL U735 ( .A(n685), .B(n43), .C(n684), .D(n25), .E(n600), .F(n19), .G(
        n601), .H(n40), .Y(n599) );
  AO2222XL U736 ( .A(n740), .B(n42), .C(n739), .D(n24), .E(n443), .F(n18), .G(
        n444), .H(n39), .Y(n442) );
  AO2222XL U737 ( .A(n725), .B(n43), .C(n724), .D(n25), .E(n503), .F(n19), .G(
        n504), .H(n40), .Y(n502) );
  AO2222XL U738 ( .A(n715), .B(n42), .C(n714), .D(n24), .E(n479), .F(n18), .G(
        n480), .H(n39), .Y(n478) );
  AO2222XL U739 ( .A(n730), .B(n42), .C(n729), .D(n24), .E(n515), .F(n18), .G(
        n516), .H(n39), .Y(n514) );
  AO2222XL U740 ( .A(n740), .B(n30), .C(n739), .D(n27), .E(n443), .F(n21), .G(
        n444), .H(n15), .Y(n449) );
  AO2222XL U741 ( .A(n715), .B(n31), .C(n714), .D(n28), .E(n479), .F(n22), .G(
        n480), .H(n16), .Y(n485) );
  AO2222XL U742 ( .A(n730), .B(n30), .C(n729), .D(n27), .E(n515), .F(n21), .G(
        n516), .H(n15), .Y(n521) );
  AO2222XL U743 ( .A(n688), .B(n31), .C(n687), .D(n28), .E(n575), .F(n22), .G(
        n576), .H(n16), .Y(n581) );
  OAI221X1 U744 ( .A(n45), .B(n553), .C(n47), .D(n554), .E(n555), .Y(n549) );
  AOI32X1 U745 ( .A(n9), .B(n695), .C(n552), .D(n551), .E(n36), .Y(n555) );
  OAI221X1 U746 ( .A(n44), .B(n553), .C(n46), .D(n554), .E(n558), .Y(n556) );
  AOI32X1 U747 ( .A(n33), .B(n695), .C(n552), .D(n551), .E(n12), .Y(n558) );
  OAI221X1 U748 ( .A(n45), .B(n529), .C(n47), .D(n530), .E(n531), .Y(n525) );
  AOI32X1 U749 ( .A(n10), .B(n238), .C(n528), .D(n527), .E(n37), .Y(n531) );
  OAI221X1 U750 ( .A(n44), .B(n529), .C(n46), .D(n530), .E(n534), .Y(n532) );
  AOI32X1 U751 ( .A(n33), .B(n238), .C(n528), .D(n527), .E(n13), .Y(n534) );
  OAI221X1 U752 ( .A(n44), .B(n619), .C(n46), .D(n620), .E(n624), .Y(n622) );
  AOI32X1 U753 ( .A(n34), .B(n673), .C(n618), .D(n617), .E(n13), .Y(n624) );
  OAI221X1 U754 ( .A(n45), .B(n619), .C(n47), .D(n620), .E(n621), .Y(n615) );
  AOI32X1 U755 ( .A(n10), .B(n673), .C(n618), .D(n617), .E(n37), .Y(n621) );
  AOI22X1 U756 ( .A(n314), .B(n80), .C(n315), .D(n80), .Y(n426) );
  INVX1 U757 ( .A(N1217), .Y(n103) );
  AO21X1 U758 ( .B(n72), .C(n150), .A(n149), .Y(n172) );
  INVX1 U759 ( .A(n665), .Y(n150) );
  MUX4X1 U760 ( .D0(n649), .D1(n648), .D2(n642), .D3(n641), .S0(n3), .S1(n76), 
        .Y(n149) );
  AO2222XL U761 ( .A(n667), .B(n42), .C(n666), .D(n24), .E(n643), .F(n18), .G(
        n644), .H(n39), .Y(n642) );
  MUX2X1 U762 ( .D0(n143), .D1(n142), .S(cs_ptr[0]), .Y(n179) );
  AO21X1 U763 ( .B(n6), .C(n141), .A(n139), .Y(n143) );
  AO21X1 U764 ( .B(n4), .C(n141), .A(n140), .Y(n142) );
  INVX1 U765 ( .A(n669), .Y(n141) );
  AO2222XL U766 ( .A(n704), .B(n43), .C(n703), .D(n25), .E(n527), .F(n19), .G(
        n528), .H(n40), .Y(n526) );
  MUX2X1 U767 ( .D0(n637), .D1(n636), .S(n57), .Y(n140) );
  AO2222XL U768 ( .A(n30), .B(n671), .C(n27), .D(n670), .E(n21), .F(n631), .G(
        n15), .H(n632), .Y(n637) );
  OAI221X1 U769 ( .A(n633), .B(n44), .C(n634), .D(n46), .E(n638), .Y(n636) );
  AOI32X1 U770 ( .A(n632), .B(n669), .C(n34), .D(n12), .E(n631), .Y(n638) );
  OAI22AX1 U771 ( .D(n76), .C(n451), .A(n78), .B(n452), .Y(n433) );
  AOI222XL U772 ( .A(N1225), .B(n4), .C(n460), .D(n733), .E(N1224), .F(n461), 
        .Y(n451) );
  AOI222XL U773 ( .A(N1225), .B(n7), .C(n453), .D(n733), .E(N1224), .F(n454), 
        .Y(n452) );
  INVX1 U774 ( .A(N1224), .Y(n733) );
  OAI221X1 U775 ( .A(n745), .B(n457), .C(n743), .D(n458), .E(n459), .Y(n453)
         );
  AOI32X1 U776 ( .A(n10), .B(n732), .C(n456), .D(n455), .E(n37), .Y(n459) );
  OAI221X1 U777 ( .A(n744), .B(n457), .C(n742), .D(n458), .E(n462), .Y(n460)
         );
  AOI32X1 U778 ( .A(n34), .B(n732), .C(n456), .D(n455), .E(n13), .Y(n462) );
  OAI221X1 U779 ( .A(n44), .B(n645), .C(n46), .D(n646), .E(n650), .Y(n648) );
  AOI32X1 U780 ( .A(n33), .B(n665), .C(n644), .D(n643), .E(n12), .Y(n650) );
  MUX2X1 U781 ( .D0(n630), .D1(n629), .S(n57), .Y(n139) );
  AO2222XL U782 ( .A(n42), .B(n671), .C(n24), .D(n670), .E(n18), .F(n631), .G(
        n39), .H(n632), .Y(n630) );
  OAI221X1 U783 ( .A(n633), .B(n45), .C(n634), .D(n47), .E(n635), .Y(n629) );
  AOI32X1 U784 ( .A(n632), .B(n669), .C(n9), .D(n36), .E(n631), .Y(n635) );
  OAI221X1 U785 ( .A(n45), .B(n645), .C(n47), .D(n646), .E(n647), .Y(n641) );
  AOI32X1 U786 ( .A(n9), .B(n665), .C(n644), .D(n643), .E(n36), .Y(n647) );
  INVX1 U787 ( .A(N1795), .Y(n81) );
  AO2222XL U788 ( .A(n698), .B(n42), .C(n697), .D(n24), .E(n551), .F(n18), .G(
        n552), .H(n39), .Y(n550) );
  AO2222XL U789 ( .A(n735), .B(n43), .C(n734), .D(n25), .E(n455), .F(n19), .G(
        n456), .H(n40), .Y(n454) );
  AO2222XL U790 ( .A(n698), .B(n30), .C(n697), .D(n27), .E(n551), .F(n21), .G(
        n552), .H(n15), .Y(n557) );
  AO2222XL U791 ( .A(n735), .B(n31), .C(n734), .D(n28), .E(n455), .F(n22), .G(
        n456), .H(n16), .Y(n461) );
  AO2222XL U792 ( .A(n667), .B(n30), .C(n666), .D(n27), .E(n643), .F(n21), .G(
        n644), .H(n15), .Y(n649) );
  INVX1 U793 ( .A(r_dac_en[7]), .Y(n742) );
  INVX1 U794 ( .A(r_dac_en[5]), .Y(n744) );
  INVX1 U795 ( .A(r_dac_en[4]), .Y(n745) );
  INVX1 U796 ( .A(r_dac_en[6]), .Y(n743) );
  INVX1 U797 ( .A(r_dac_en[17]), .Y(n245) );
  NOR2X1 U798 ( .A(pos_dacis[9]), .B(pos_dacis[8]), .Y(n289) );
  NAND4X1 U799 ( .A(n757), .B(n758), .C(n288), .D(n759), .Y(n286) );
  NOR2X1 U800 ( .A(pos_dacis[17]), .B(pos_dacis[16]), .Y(n288) );
  INVX1 U801 ( .A(r_comp_swtch), .Y(n365) );
  INVXL U802 ( .A(n230), .Y(n223) );
  NAND32XL U803 ( .B(n219), .C(n218), .A(n217), .Y(n230) );
  OAI211X1 U804 ( .C(n186), .D(n383), .A(n185), .B(n184), .Y(n760) );
  AND2XL U805 ( .A(n391), .B(ps_ptr[4]), .Y(N1035) );
  INVXL U806 ( .A(ps_ptr[4]), .Y(n297) );
  INVX4 U807 ( .A(n153), .Y(n180) );
  AOI31X1 U808 ( .A(n398), .B(n399), .C(n397), .D(n281), .Y(n215) );
  NAND21X2 U809 ( .B(n172), .A(n178), .Y(n153) );
  AND3X2 U810 ( .A(n235), .B(n234), .C(n233), .Y(n242) );
  OA222X1 U811 ( .A(n183), .B(n271), .C(n182), .D(n218), .E(n181), .F(n274), 
        .Y(n184) );
  NAND21XL U812 ( .B(ps_ptr[4]), .A(n320), .Y(n321) );
  OAI22XL U813 ( .A(ps_ptr[4]), .B(n103), .C(ps_ptr[3]), .D(n99), .Y(n295) );
  AOI211X1 U814 ( .C(n232), .D(n103), .A(n231), .B(n230), .Y(n233) );
  NAND21X4 U815 ( .B(r_semi), .A(n151), .Y(n152) );
  NAND32X4 U816 ( .B(n179), .C(n155), .A(n180), .Y(n275) );
  XNOR2XL U817 ( .A(N1586), .B(sub_395_S2_I11_aco_carry[5]), .Y(N1595) );
  XNOR2XL U818 ( .A(N1504), .B(sub_395_S2_I9_aco_carry[5]), .Y(N1513) );
  XNOR2XL U819 ( .A(N1709), .B(sub_395_S2_I14_aco_carry[5]), .Y(N1718) );
  XNOR2XL U820 ( .A(N1463), .B(sub_395_S2_I8_aco_carry[5]), .Y(N1472) );
  XNOR2XL U821 ( .A(N1299), .B(sub_395_S2_I4_aco_carry[5]), .Y(N1308) );
  XNOR2XL U822 ( .A(n102), .B(sub_395_S2_I2_aco_carry[5]), .Y(N1226) );
  XNOR2XL U823 ( .A(N1422), .B(sub_395_S2_I7_aco_carry[5]), .Y(N1431) );
  XNOR2XL U824 ( .A(N1258), .B(sub_395_S2_I3_aco_carry[5]), .Y(N1267) );
  XNOR2XL U825 ( .A(N1381), .B(sub_395_S2_I6_aco_carry[5]), .Y(N1390) );
  XNOR2XL U826 ( .A(N1340), .B(sub_395_S2_I5_aco_carry[5]), .Y(N1349) );
  XNOR2XL U827 ( .A(N1176), .B(sub_395_S2_aco_carry[5]), .Y(N1185) );
  XNOR2XL U828 ( .A(N1668), .B(sub_395_S2_I13_aco_carry[5]), .Y(N1677) );
  XNOR2XL U829 ( .A(N1627), .B(sub_395_S2_I12_aco_carry[5]), .Y(N1636) );
  OR2X1 U830 ( .A(sub_395_S2_aco_carry[3]), .B(N1174), .Y(
        sub_395_S2_aco_carry[4]) );
  XNOR2XL U831 ( .A(sub_395_S2_aco_carry[3]), .B(N1174), .Y(N1183) );
  OR2X1 U832 ( .A(sub_395_S2_aco_carry[2]), .B(N1173), .Y(
        sub_395_S2_aco_carry[3]) );
  XNOR2XL U833 ( .A(sub_395_S2_aco_carry[2]), .B(N1173), .Y(N1182) );
  OR2X1 U834 ( .A(N1172), .B(n55), .Y(sub_395_S2_aco_carry[2]) );
  XNOR2XL U835 ( .A(N1172), .B(n55), .Y(N1181) );
  OR2X1 U836 ( .A(add_394_carry_4_), .B(N1217), .Y(N1176) );
  XNOR2XL U837 ( .A(add_394_carry_4_), .B(N1217), .Y(N1175) );
  AND2X1 U838 ( .A(n95), .B(add_394_carry_3_), .Y(add_394_carry_4_) );
  XOR2X1 U839 ( .A(add_394_carry_3_), .B(n95), .Y(N1174) );
  AND2X1 U840 ( .A(n89), .B(add_394_carry_2_), .Y(add_394_carry_3_) );
  XOR2X1 U841 ( .A(add_394_carry_2_), .B(cs_ptr[2]), .Y(N1173) );
  AND2X1 U842 ( .A(n83), .B(n76), .Y(add_394_carry_2_) );
  XOR2X1 U843 ( .A(cs_ptr[0]), .B(cs_ptr[1]), .Y(N1172) );
  OR2X1 U844 ( .A(sub_395_S2_I2_aco_carry[3]), .B(n97), .Y(
        sub_395_S2_I2_aco_carry[4]) );
  XNOR2XL U845 ( .A(sub_395_S2_I2_aco_carry[3]), .B(n96), .Y(N1224) );
  OR2X1 U846 ( .A(sub_395_S2_I2_aco_carry[2]), .B(n91), .Y(
        sub_395_S2_I2_aco_carry[3]) );
  XNOR2XL U847 ( .A(sub_395_S2_I2_aco_carry[2]), .B(n90), .Y(N1223) );
  OR2X1 U848 ( .A(N1705), .B(n71), .Y(sub_395_S2_I2_aco_carry[2]) );
  XNOR2XL U849 ( .A(n84), .B(n71), .Y(N1222) );
  OR2X1 U850 ( .A(sub_395_S2_I5_aco_carry[3]), .B(N1338), .Y(
        sub_395_S2_I5_aco_carry[4]) );
  XNOR2XL U851 ( .A(sub_395_S2_I5_aco_carry[3]), .B(N1338), .Y(N1347) );
  OR2X1 U852 ( .A(sub_395_S2_I5_aco_carry[2]), .B(N1337), .Y(
        sub_395_S2_I5_aco_carry[3]) );
  XNOR2XL U853 ( .A(sub_395_S2_I5_aco_carry[2]), .B(N1337), .Y(N1346) );
  OR2X1 U854 ( .A(N1336), .B(n54), .Y(sub_395_S2_I5_aco_carry[2]) );
  XNOR2XL U855 ( .A(N1336), .B(n54), .Y(N1345) );
  AND2X1 U856 ( .A(n102), .B(add_394_I5_carry_4_), .Y(N1340) );
  XOR2X1 U857 ( .A(add_394_I5_carry_4_), .B(n101), .Y(N1339) );
  OR2X1 U858 ( .A(add_394_I5_carry_3_), .B(n97), .Y(add_394_I5_carry_4_) );
  XNOR2XL U859 ( .A(add_394_I5_carry_3_), .B(n97), .Y(N1338) );
  OR2X1 U860 ( .A(add_394_I5_carry_2_), .B(n91), .Y(add_394_I5_carry_3_) );
  XNOR2XL U861 ( .A(add_394_I5_carry_2_), .B(n90), .Y(N1337) );
  AND2X1 U862 ( .A(n83), .B(n76), .Y(add_394_I5_carry_2_) );
  XOR2X1 U863 ( .A(cs_ptr[0]), .B(cs_ptr[1]), .Y(N1336) );
  OR2X1 U864 ( .A(sub_395_S2_I6_aco_carry[3]), .B(N1379), .Y(
        sub_395_S2_I6_aco_carry[4]) );
  XNOR2XL U865 ( .A(sub_395_S2_I6_aco_carry[3]), .B(N1379), .Y(N1388) );
  OR2X1 U866 ( .A(sub_395_S2_I6_aco_carry[2]), .B(n92), .Y(
        sub_395_S2_I6_aco_carry[3]) );
  XNOR2XL U867 ( .A(sub_395_S2_I6_aco_carry[2]), .B(n93), .Y(N1387) );
  OR2X1 U868 ( .A(cs_ptr[1]), .B(n68), .Y(sub_395_S2_I6_aco_carry[2]) );
  XNOR2XL U869 ( .A(n84), .B(n68), .Y(N1386) );
  AND2X1 U870 ( .A(n101), .B(add_394_I6_carry_4_), .Y(N1381) );
  XOR2X1 U871 ( .A(add_394_I6_carry_4_), .B(n101), .Y(N1380) );
  OR2X1 U872 ( .A(cs_ptr[2]), .B(n96), .Y(add_394_I6_carry_4_) );
  XNOR2XL U873 ( .A(n89), .B(n96), .Y(N1379) );
  OR2X1 U874 ( .A(sub_395_S2_I7_aco_carry[3]), .B(N1420), .Y(
        sub_395_S2_I7_aco_carry[4]) );
  XNOR2XL U875 ( .A(sub_395_S2_I7_aco_carry[3]), .B(N1420), .Y(N1429) );
  OR2X1 U876 ( .A(sub_395_S2_I7_aco_carry[2]), .B(N1419), .Y(
        sub_395_S2_I7_aco_carry[3]) );
  XNOR2XL U877 ( .A(sub_395_S2_I7_aco_carry[2]), .B(N1419), .Y(N1428) );
  OR2X1 U878 ( .A(N1418), .B(n52), .Y(sub_395_S2_I7_aco_carry[2]) );
  XNOR2XL U879 ( .A(N1418), .B(n52), .Y(N1427) );
  AND2X1 U880 ( .A(n101), .B(add_394_I7_carry_4_), .Y(N1422) );
  XOR2X1 U881 ( .A(add_394_I7_carry_4_), .B(n101), .Y(N1421) );
  OR2X1 U882 ( .A(add_394_I7_carry_3_), .B(n97), .Y(add_394_I7_carry_4_) );
  XNOR2XL U883 ( .A(add_394_I7_carry_3_), .B(n97), .Y(N1420) );
  AND2X1 U884 ( .A(n89), .B(add_394_I7_carry_2_), .Y(add_394_I7_carry_3_) );
  XOR2X1 U885 ( .A(add_394_I7_carry_2_), .B(cs_ptr[2]), .Y(N1419) );
  OR2X1 U886 ( .A(n77), .B(n85), .Y(add_394_I7_carry_2_) );
  XNOR2XL U887 ( .A(n76), .B(n85), .Y(N1418) );
  OR2X1 U888 ( .A(sub_395_S2_I4_aco_carry[3]), .B(N1297), .Y(
        sub_395_S2_I4_aco_carry[4]) );
  XNOR2XL U889 ( .A(sub_395_S2_I4_aco_carry[3]), .B(N1297), .Y(N1306) );
  OR2X1 U890 ( .A(sub_395_S2_I4_aco_carry[2]), .B(N1296), .Y(
        sub_395_S2_I4_aco_carry[3]) );
  XNOR2XL U891 ( .A(sub_395_S2_I4_aco_carry[2]), .B(N1296), .Y(N1305) );
  OR2X1 U892 ( .A(n86), .B(n67), .Y(sub_395_S2_I4_aco_carry[2]) );
  XNOR2XL U893 ( .A(n87), .B(n67), .Y(N1304) );
  AND2X1 U894 ( .A(n101), .B(add_394_I4_carry[4]), .Y(N1299) );
  XOR2X1 U895 ( .A(add_394_I4_carry[4]), .B(n101), .Y(N1298) );
  OR2X1 U896 ( .A(add_394_I4_carry[3]), .B(n96), .Y(add_394_I4_carry[4]) );
  XNOR2XL U897 ( .A(add_394_I4_carry[3]), .B(cs_ptr[3]), .Y(N1297) );
  OR2X1 U898 ( .A(n85), .B(n91), .Y(add_394_I4_carry[3]) );
  XNOR2XL U899 ( .A(n84), .B(n90), .Y(N1296) );
  OR2X1 U900 ( .A(sub_395_S2_I3_aco_carry[3]), .B(N1256), .Y(
        sub_395_S2_I3_aco_carry[4]) );
  XNOR2XL U901 ( .A(sub_395_S2_I3_aco_carry[3]), .B(N1256), .Y(N1265) );
  OR2X1 U902 ( .A(sub_395_S2_I3_aco_carry[2]), .B(N1255), .Y(
        sub_395_S2_I3_aco_carry[3]) );
  XNOR2XL U903 ( .A(sub_395_S2_I3_aco_carry[2]), .B(N1255), .Y(N1264) );
  OR2X1 U904 ( .A(N1254), .B(n56), .Y(sub_395_S2_I3_aco_carry[2]) );
  XNOR2XL U905 ( .A(N1254), .B(n56), .Y(N1263) );
  AND2X1 U906 ( .A(n101), .B(add_394_I3_carry_4_), .Y(N1258) );
  XOR2X1 U907 ( .A(add_394_I3_carry_4_), .B(n101), .Y(N1257) );
  OR2X1 U908 ( .A(add_394_I3_carry_3_), .B(n96), .Y(add_394_I3_carry_4_) );
  XNOR2XL U909 ( .A(add_394_I3_carry_3_), .B(n97), .Y(N1256) );
  OR2X1 U910 ( .A(add_394_I3_carry_2_), .B(n91), .Y(add_394_I3_carry_3_) );
  XNOR2XL U911 ( .A(add_394_I3_carry_2_), .B(n90), .Y(N1255) );
  OR2X1 U912 ( .A(n77), .B(n85), .Y(add_394_I3_carry_2_) );
  XNOR2XL U913 ( .A(n76), .B(n85), .Y(N1254) );
  OR2X1 U914 ( .A(sub_395_S2_I8_aco_carry[3]), .B(N1461), .Y(
        sub_395_S2_I8_aco_carry[4]) );
  OR2X1 U915 ( .A(sub_395_S2_I8_aco_carry[2]), .B(N1460), .Y(
        sub_395_S2_I8_aco_carry[3]) );
  OR2X1 U916 ( .A(n86), .B(n413), .Y(sub_395_S2_I8_aco_carry[2]) );
  AND2X1 U917 ( .A(n101), .B(add_394_I8_carry[4]), .Y(N1463) );
  XOR2X1 U918 ( .A(add_394_I8_carry[4]), .B(cs_ptr[4]), .Y(N1462) );
  OR2X1 U919 ( .A(add_394_I8_carry[3]), .B(n96), .Y(add_394_I8_carry[4]) );
  XNOR2XL U920 ( .A(add_394_I8_carry[3]), .B(n97), .Y(N1461) );
  AND2X1 U921 ( .A(n89), .B(n83), .Y(add_394_I8_carry[3]) );
  XOR2X1 U922 ( .A(cs_ptr[1]), .B(cs_ptr[2]), .Y(N1460) );
  OR2X1 U923 ( .A(sub_395_S2_I9_aco_carry[3]), .B(N1502), .Y(
        sub_395_S2_I9_aco_carry[4]) );
  OR2X1 U924 ( .A(sub_395_S2_I9_aco_carry[2]), .B(N1501), .Y(
        sub_395_S2_I9_aco_carry[3]) );
  OR2X1 U925 ( .A(N1500), .B(n414), .Y(sub_395_S2_I9_aco_carry[2]) );
  AND2X1 U926 ( .A(n102), .B(add_394_I9_carry_4_), .Y(N1504) );
  XOR2X1 U927 ( .A(add_394_I9_carry_4_), .B(cs_ptr[4]), .Y(N1503) );
  OR2X1 U928 ( .A(add_394_I9_carry_3_), .B(n96), .Y(add_394_I9_carry_4_) );
  XNOR2XL U929 ( .A(add_394_I9_carry_3_), .B(n97), .Y(N1502) );
  AND2X1 U930 ( .A(n89), .B(add_394_I9_carry_2_), .Y(add_394_I9_carry_3_) );
  XOR2X1 U931 ( .A(add_394_I9_carry_2_), .B(cs_ptr[2]), .Y(N1501) );
  AND2X1 U932 ( .A(n83), .B(n76), .Y(add_394_I9_carry_2_) );
  XOR2X1 U933 ( .A(cs_ptr[0]), .B(cs_ptr[1]), .Y(N1500) );
  OR2X1 U934 ( .A(sub_395_S2_I10_aco_carry[3]), .B(n98), .Y(
        sub_395_S2_I10_aco_carry[4]) );
  OR2X1 U935 ( .A(sub_395_S2_I10_aco_carry[2]), .B(n91), .Y(
        sub_395_S2_I10_aco_carry[3]) );
  OR2X1 U936 ( .A(N1705), .B(n415), .Y(sub_395_S2_I10_aco_carry[2]) );
  AND2X1 U937 ( .A(n102), .B(n97), .Y(N1545) );
  XOR2X1 U938 ( .A(cs_ptr[3]), .B(cs_ptr[4]), .Y(N1544) );
  OR2X1 U939 ( .A(sub_395_S2_I11_aco_carry[3]), .B(N1584), .Y(
        sub_395_S2_I11_aco_carry[4]) );
  XNOR2XL U940 ( .A(sub_395_S2_I11_aco_carry[3]), .B(N1584), .Y(N1593) );
  OR2X1 U941 ( .A(sub_395_S2_I11_aco_carry[2]), .B(N1583), .Y(
        sub_395_S2_I11_aco_carry[3]) );
  XNOR2XL U942 ( .A(sub_395_S2_I11_aco_carry[2]), .B(N1583), .Y(N1592) );
  OR2X1 U943 ( .A(N1582), .B(n53), .Y(sub_395_S2_I11_aco_carry[2]) );
  XNOR2XL U944 ( .A(N1582), .B(n53), .Y(N1591) );
  AND2X1 U945 ( .A(n102), .B(add_394_I11_carry_4_), .Y(N1586) );
  XOR2X1 U946 ( .A(add_394_I11_carry_4_), .B(cs_ptr[4]), .Y(N1585) );
  AND2X1 U947 ( .A(n97), .B(add_394_I11_carry_3_), .Y(add_394_I11_carry_4_) );
  XOR2X1 U948 ( .A(add_394_I11_carry_3_), .B(n95), .Y(N1584) );
  OR2X1 U949 ( .A(add_394_I11_carry_2_), .B(n91), .Y(add_394_I11_carry_3_) );
  XNOR2XL U950 ( .A(add_394_I11_carry_2_), .B(n90), .Y(N1583) );
  OR2X1 U951 ( .A(n78), .B(n85), .Y(add_394_I11_carry_2_) );
  XNOR2XL U952 ( .A(n76), .B(n85), .Y(N1582) );
  OR2X1 U953 ( .A(sub_395_S2_I12_aco_carry[3]), .B(N1625), .Y(
        sub_395_S2_I12_aco_carry[4]) );
  OR2X1 U954 ( .A(sub_395_S2_I12_aco_carry[2]), .B(N1624), .Y(
        sub_395_S2_I12_aco_carry[3]) );
  OR2X1 U955 ( .A(n86), .B(n416), .Y(sub_395_S2_I12_aco_carry[2]) );
  AND2X1 U956 ( .A(n102), .B(add_394_I12_carry[4]), .Y(N1627) );
  XOR2X1 U957 ( .A(add_394_I12_carry[4]), .B(cs_ptr[4]), .Y(N1626) );
  AND2X1 U958 ( .A(n95), .B(add_394_I12_carry[3]), .Y(add_394_I12_carry[4]) );
  XOR2X1 U959 ( .A(add_394_I12_carry[3]), .B(n95), .Y(N1625) );
  OR2X1 U960 ( .A(cs_ptr[1]), .B(n91), .Y(add_394_I12_carry[3]) );
  XNOR2XL U961 ( .A(n84), .B(n90), .Y(N1624) );
  OR2X1 U962 ( .A(sub_395_S2_I14_aco_carry[3]), .B(N1707), .Y(
        sub_395_S2_I14_aco_carry[4]) );
  XNOR2XL U963 ( .A(sub_395_S2_I14_aco_carry[3]), .B(N1707), .Y(N1716) );
  OR2X1 U964 ( .A(sub_395_S2_I14_aco_carry[2]), .B(n92), .Y(
        sub_395_S2_I14_aco_carry[3]) );
  XNOR2XL U965 ( .A(sub_395_S2_I14_aco_carry[2]), .B(n92), .Y(N1715) );
  OR2X1 U966 ( .A(cs_ptr[1]), .B(n66), .Y(sub_395_S2_I14_aco_carry[2]) );
  XNOR2XL U967 ( .A(n84), .B(n66), .Y(N1714) );
  AND2X1 U968 ( .A(n102), .B(add_394_I14_carry_4_), .Y(N1709) );
  XOR2X1 U969 ( .A(add_394_I14_carry_4_), .B(cs_ptr[4]), .Y(N1708) );
  AND2X1 U970 ( .A(n95), .B(n89), .Y(add_394_I14_carry_4_) );
  XOR2X1 U971 ( .A(cs_ptr[2]), .B(cs_ptr[3]), .Y(N1707) );
  OR2X1 U972 ( .A(sub_395_S2_I13_aco_carry[3]), .B(N1666), .Y(
        sub_395_S2_I13_aco_carry[4]) );
  OR2X1 U973 ( .A(sub_395_S2_I13_aco_carry[2]), .B(N1665), .Y(
        sub_395_S2_I13_aco_carry[3]) );
  OR2X1 U974 ( .A(N1664), .B(n417), .Y(sub_395_S2_I13_aco_carry[2]) );
  AND2X1 U975 ( .A(n102), .B(add_394_I13_carry_4_), .Y(N1668) );
  XOR2X1 U976 ( .A(add_394_I13_carry_4_), .B(cs_ptr[4]), .Y(N1667) );
  AND2X1 U977 ( .A(n95), .B(add_394_I13_carry_3_), .Y(add_394_I13_carry_4_) );
  XOR2X1 U978 ( .A(add_394_I13_carry_3_), .B(cs_ptr[3]), .Y(N1666) );
  OR2X1 U979 ( .A(add_394_I13_carry_2_), .B(n91), .Y(add_394_I13_carry_3_) );
  XNOR2XL U980 ( .A(add_394_I13_carry_2_), .B(n90), .Y(N1665) );
  AND2X1 U981 ( .A(n83), .B(n76), .Y(add_394_I13_carry_2_) );
  XOR2X1 U982 ( .A(cs_ptr[0]), .B(cs_ptr[1]), .Y(N1664) );
  AND2X1 U983 ( .A(n102), .B(add_394_I15_carry_4_), .Y(N1750) );
  AND2X1 U984 ( .A(n95), .B(add_394_I15_carry_3_), .Y(add_394_I15_carry_4_) );
  AND2X1 U985 ( .A(n89), .B(add_394_I15_carry_2_), .Y(add_394_I15_carry_3_) );
  OR2X1 U986 ( .A(n78), .B(n85), .Y(add_394_I15_carry_2_) );
  AND2X1 U987 ( .A(n95), .B(add_394_I16_carry[3]), .Y(add_394_I16_carry[4]) );
  AND2X1 U988 ( .A(n89), .B(n83), .Y(add_394_I16_carry[3]) );
  AOI21X1 U989 ( .B(N1708), .C(N1707), .A(N1709), .Y(n425) );
  OAI21X1 U990 ( .B(n93), .C(n84), .A(N1708), .Y(n418) );
  AOI21X1 U991 ( .B(N1667), .C(N1666), .A(N1668), .Y(n609) );
  OAI21X1 U992 ( .B(N1665), .C(N1664), .A(N1667), .Y(n608) );
  NAND2X1 U993 ( .A(n609), .B(n608), .Y(N1669) );
  AOI21X1 U994 ( .B(N1626), .C(N1625), .A(N1627), .Y(n611) );
  OAI21X1 U995 ( .B(N1624), .C(n86), .A(N1626), .Y(n610) );
  NAND2X1 U996 ( .A(n611), .B(n610), .Y(N1628) );
  AOI21X1 U997 ( .B(N1585), .C(N1584), .A(N1586), .Y(n613) );
  OAI21X1 U998 ( .B(N1583), .C(N1582), .A(N1585), .Y(n612) );
  AOI21X1 U999 ( .B(N1544), .C(n98), .A(N1545), .Y(n625) );
  OAI21X1 U1000 ( .B(n89), .C(n84), .A(N1544), .Y(n614) );
  NAND2X1 U1001 ( .A(n625), .B(n614), .Y(N1546) );
  AOI21X1 U1002 ( .B(N1503), .C(N1502), .A(N1504), .Y(n627) );
  OAI21X1 U1003 ( .B(N1501), .C(N1500), .A(N1503), .Y(n626) );
  NAND2X1 U1004 ( .A(n627), .B(n626), .Y(N1505) );
  AOI21X1 U1005 ( .B(N1462), .C(N1461), .A(N1463), .Y(n639) );
  OAI21X1 U1006 ( .B(N1460), .C(n86), .A(N1462), .Y(n628) );
  NAND2X1 U1007 ( .A(n639), .B(n628), .Y(N1464) );
  AOI21X1 U1008 ( .B(N1421), .C(N1420), .A(N1422), .Y(n651) );
  OAI21X1 U1009 ( .B(N1419), .C(N1418), .A(N1421), .Y(n640) );
  AOI21X1 U1010 ( .B(N1380), .C(N1379), .A(N1381), .Y(n653) );
  OAI21X1 U1011 ( .B(n92), .C(n84), .A(N1380), .Y(n652) );
  AOI21X1 U1012 ( .B(N1339), .C(N1338), .A(N1340), .Y(n655) );
  OAI21X1 U1013 ( .B(N1337), .C(N1336), .A(N1339), .Y(n654) );
  AOI21X1 U1014 ( .B(N1298), .C(N1297), .A(N1299), .Y(n657) );
  OAI21X1 U1015 ( .B(N1296), .C(n86), .A(N1298), .Y(n656) );
  AOI21X1 U1016 ( .B(N1257), .C(N1256), .A(N1258), .Y(n659) );
  OAI21X1 U1017 ( .B(N1255), .C(N1254), .A(N1257), .Y(n658) );
  AOI21X1 U1018 ( .B(n103), .C(n96), .A(n102), .Y(n662) );
  OAI21X1 U1019 ( .B(n90), .C(n84), .A(n104), .Y(n661) );
  AOI21X1 U1020 ( .B(N1175), .C(N1174), .A(N1176), .Y(n664) );
  OAI21X1 U1021 ( .B(N1173), .C(N1172), .A(N1175), .Y(n663) );
endmodule


module SNPS_CLOCK_GATE_HIGH_shmux_00000005_00000012_00000012_1 ( CLK, EN, 
        ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_shmux_00000005_00000012_00000012_0 ( CLK, EN, 
        ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module dac2sar_a0 ( r_dac_t, r_dacyc, r_sar10, sar_ini, sar_nxt, semi_nxt, 
        auto_sar, busy, stop, sync_i, sampl_begn, sampl_done, sh_rst, 
        dacyc_done, sacyc_done, dac_v, rpt_v, clk, srstz );
  input [1:0] r_dac_t;
  output [9:0] dac_v;
  output [9:0] rpt_v;
  input r_dacyc, r_sar10, sar_ini, sar_nxt, semi_nxt, auto_sar, busy, stop,
         sync_i, clk, srstz;
  output sampl_begn, sampl_done, sh_rst, dacyc_done, sacyc_done;
  wire   n124, N19, N20, N21, N23, N36, N37, N38, N39, N40, N41, N42, N43, N44,
         N45, N46, N47, N48, N49, N50, N60, N61, N62, N63, N64, N68, updlo,
         updup, upd1v, N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N82,
         N83, N84, N85, N86, N87, N88, N89, N90, N91, net10186, net10192, n55,
         n56, n57, n58, n61, n62, n63, n64, n65, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n97, n98, n103, n104, n105, n106, n107,
         n108, n109, n4, n5, n6, n7, n8, n9, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n59, n60, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n99, n100, n101, n102, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123,
         SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2,
         SYNOPSYS_UNCONNECTED_3;
  wire   [6:0] dacnt;
  wire   [3:0] sarcyc;
  wire   [9:0] r_lt_lo;
  wire   [9:0] r_lt_up;
  wire   [9:0] r_avg00;
  wire   [9:0] r_avgup;
  wire   [9:0] r_dacvo;

  glreg_WIDTH10_2 u0_dac1v ( .clk(clk), .arstz(n26), .we(upd1v), .wdat(r_dacvo), .rdat({dac_v[9:1], n124}) );
  glreg_WIDTH10_1 u0_lt_lo ( .clk(clk), .arstz(n25), .we(updlo), .wdat({n6, n4, 
        n15, n5, n17, n16, n13, n12, n14, n18}), .rdat(r_lt_lo) );
  glreg_WIDTH10_0 u0_lt_up ( .clk(clk), .arstz(n24), .we(updup), .wdat(r_avgup), .rdat(r_lt_up) );
  SNPS_CLOCK_GATE_HIGH_dac2sar_a0_0 clk_gate_dacnt_reg ( .CLK(clk), .EN(N43), 
        .ENCLK(net10186), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_dac2sar_a0_1 clk_gate_sarcyc_reg ( .CLK(clk), .EN(N60), 
        .ENCLK(net10192), .TE(1'b0) );
  dac2sar_a0_DW01_add_0 add_303 ( .A({1'b0, n96, n99, n101, n110, n112, n114, 
        n116, n118, n120, n122}), .B({1'b0, n95, n100, n102, n111, n113, n115, 
        n117, n119, n121, n123}), .CI(1'b0), .SUM({N91, N90, N89, N88, N87, 
        N86, N85, N84, N83, N82, SYNOPSYS_UNCONNECTED_1}), .CO() );
  dac2sar_a0_DW01_add_2 add_296 ( .A({1'b0, r_lt_lo}), .B({1'b0, r_lt_up}), 
        .CI(1'b0), .SUM({r_avg00, SYNOPSYS_UNCONNECTED_2}), .CO() );
  dac2sar_a0_DW01_inc_0 add_276 ( .A(dacnt), .SUM({N42, N41, N40, N39, N38, 
        N37, N36}) );
  dac2sar_a0_DW01_add_3 add_301 ( .A({1'b0, n6, n4, n15, n5, n17, n16, n13, 
        n12, n14, n18}), .B({1'b0, r_avgup}), .CI(1'b0), .SUM({N80, N79, N78, 
        N77, N76, N75, N74, N73, N72, N71, SYNOPSYS_UNCONNECTED_3}), .CO() );
  DFFQX1 sarcyc_reg_2_ ( .D(N63), .C(net10192), .Q(sarcyc[2]) );
  DFFQX1 sarcyc_reg_1_ ( .D(N62), .C(net10192), .Q(sarcyc[1]) );
  DFFNQX1 sh_rst_n_reg ( .D(N68), .XC(clk), .Q(sh_rst) );
  DFFQX1 sarcyc_reg_0_ ( .D(N61), .C(net10192), .Q(sarcyc[0]) );
  DFFQX1 sarcyc_reg_3_ ( .D(N64), .C(net10192), .Q(sarcyc[3]) );
  DFFQX1 dacnt_reg_1_ ( .D(N45), .C(net10186), .Q(dacnt[1]) );
  DFFQX1 dacnt_reg_4_ ( .D(N48), .C(net10186), .Q(dacnt[4]) );
  DFFQX1 dacnt_reg_0_ ( .D(N44), .C(net10186), .Q(dacnt[0]) );
  DFFQX1 dacnt_reg_5_ ( .D(N49), .C(net10186), .Q(dacnt[5]) );
  DFFQX1 dacnt_reg_2_ ( .D(N46), .C(net10186), .Q(dacnt[2]) );
  DFFQX1 dacnt_reg_3_ ( .D(N47), .C(net10186), .Q(dacnt[3]) );
  DFFQX1 dacnt_reg_6_ ( .D(N50), .C(net10186), .Q(dacnt[6]) );
  NAND21X1 U3 ( .B(n102), .A(n37), .Y(r_avgup[7]) );
  NAND21X1 U4 ( .B(n95), .A(n37), .Y(r_avgup[9]) );
  NAND2X1 U5 ( .A(n70), .B(n37), .Y(r_avgup[0]) );
  NAND21X1 U6 ( .B(n117), .A(n37), .Y(r_avgup[3]) );
  MUX2X1 U7 ( .D0(N77), .D1(r_avg00[6]), .S(n7), .Y(r_dacvo[6]) );
  MUX2X1 U8 ( .D0(N80), .D1(r_avg00[9]), .S(semi_nxt), .Y(r_dacvo[9]) );
  MUX2X1 U9 ( .D0(N78), .D1(r_avg00[7]), .S(semi_nxt), .Y(r_dacvo[7]) );
  NOR2X1 U13 ( .A(n8), .B(n77), .Y(n4) );
  NOR2X1 U14 ( .A(sar_ini), .B(n79), .Y(n5) );
  NOR2X1 U15 ( .A(n8), .B(n76), .Y(n6) );
  BUFX3 U16 ( .A(semi_nxt), .Y(n7) );
  MUX2X1 U17 ( .D0(N76), .D1(r_avg00[5]), .S(semi_nxt), .Y(r_dacvo[5]) );
  MUX2X1 U18 ( .D0(N75), .D1(r_avg00[4]), .S(semi_nxt), .Y(r_dacvo[4]) );
  BUFX3 U19 ( .A(sar_ini), .Y(n8) );
  INVX3 U20 ( .A(sar_ini), .Y(n37) );
  INVX1 U21 ( .A(n124), .Y(n9) );
  INVX1 U22 ( .A(n9), .Y(dac_v[0]) );
  INVX1 U23 ( .A(n9), .Y(n11) );
  NAND2XL U24 ( .A(n88), .B(n37), .Y(r_avgup[6]) );
  NOR2XL U25 ( .A(sar_ini), .B(n82), .Y(n13) );
  NOR2XL U26 ( .A(sar_ini), .B(n83), .Y(n12) );
  NOR2XL U27 ( .A(sar_ini), .B(n84), .Y(n14) );
  MUX2X2 U28 ( .D0(N79), .D1(r_avg00[8]), .S(n7), .Y(r_dacvo[8]) );
  NAND2X1 U29 ( .A(n72), .B(n37), .Y(r_avgup[2]) );
  NAND21XL U30 ( .B(n113), .A(n37), .Y(r_avgup[5]) );
  NAND2XL U31 ( .A(n74), .B(n37), .Y(r_avgup[4]) );
  NOR4XL U32 ( .A(sarcyc[0]), .B(sarcyc[1]), .C(sarcyc[2]), .D(sarcyc[3]), .Y(
        n86) );
  INVX1 U33 ( .A(n27), .Y(n25) );
  INVX1 U34 ( .A(n27), .Y(n26) );
  INVX1 U35 ( .A(srstz), .Y(n27) );
  INVX1 U36 ( .A(n27), .Y(n24) );
  OR2XL U37 ( .A(stop), .B(n27), .Y(n36) );
  OR3XL U38 ( .A(sar_nxt), .B(n8), .C(semi_nxt), .Y(upd1v) );
  NAND32X1 U39 ( .B(dacyc_done), .C(n36), .A(n48), .Y(N43) );
  OR2X1 U40 ( .A(n69), .B(n34), .Y(N60) );
  INVX1 U41 ( .A(n48), .Y(n49) );
  INVX1 U42 ( .A(n53), .Y(n69) );
  INVX1 U43 ( .A(n60), .Y(n67) );
  INVX1 U44 ( .A(N23), .Y(n93) );
  MUX2X1 U45 ( .D0(N71), .D1(r_avg00[0]), .S(semi_nxt), .Y(r_dacvo[0]) );
  NAND2XL U46 ( .A(n90), .B(n37), .Y(r_avgup[8]) );
  NAND2X4 U47 ( .A(n71), .B(n37), .Y(r_avgup[1]) );
  MUX2X1 U48 ( .D0(N72), .D1(r_avg00[1]), .S(semi_nxt), .Y(r_dacvo[1]) );
  MUX2X1 U49 ( .D0(N74), .D1(r_avg00[3]), .S(semi_nxt), .Y(r_dacvo[3]) );
  MUX2X1 U50 ( .D0(N73), .D1(r_avg00[2]), .S(semi_nxt), .Y(r_dacvo[2]) );
  NOR2XL U51 ( .A(sar_ini), .B(n78), .Y(n15) );
  NOR2XL U52 ( .A(sar_ini), .B(n81), .Y(n16) );
  NOR2XL U53 ( .A(sar_ini), .B(n80), .Y(n17) );
  NOR2XL U54 ( .A(sar_ini), .B(n85), .Y(n18) );
  AO21XL U55 ( .B(sar_nxt), .C(sync_i), .A(n8), .Y(updlo) );
  NOR2X1 U56 ( .A(n92), .B(n64), .Y(sampl_begn) );
  NAND31X1 U57 ( .C(n36), .A(busy), .B(n35), .Y(n48) );
  NAND21X1 U58 ( .B(sacyc_done), .A(n33), .Y(n34) );
  INVX1 U59 ( .A(n36), .Y(n33) );
  NAND21X1 U60 ( .B(n59), .A(n69), .Y(n60) );
  NAND32X1 U61 ( .B(n35), .C(n34), .A(auto_sar), .Y(n53) );
  AND2X1 U62 ( .A(N41), .B(n49), .Y(N49) );
  AND2X1 U63 ( .A(N40), .B(n49), .Y(N48) );
  AND2X1 U64 ( .A(N39), .B(n49), .Y(N47) );
  AND2X1 U65 ( .A(N38), .B(n49), .Y(N46) );
  AND2X1 U66 ( .A(N37), .B(n49), .Y(N45) );
  AND2X1 U67 ( .A(n69), .B(n68), .Y(N61) );
  NOR2X1 U68 ( .A(N20), .B(n107), .Y(N23) );
  NOR32XL U69 ( .B(busy), .C(n92), .A(n64), .Y(N68) );
  INVX1 U70 ( .A(n90), .Y(n100) );
  INVX1 U71 ( .A(n77), .Y(n99) );
  INVX1 U72 ( .A(n76), .Y(n96) );
  INVX1 U73 ( .A(n91), .Y(n95) );
  INVX1 U74 ( .A(r_avg00[8]), .Y(n39) );
  INVX1 U75 ( .A(n83), .Y(n118) );
  INVX1 U76 ( .A(n72), .Y(n119) );
  INVX1 U77 ( .A(n82), .Y(n116) );
  INVX1 U78 ( .A(n73), .Y(n117) );
  INVX1 U79 ( .A(n81), .Y(n114) );
  INVX1 U80 ( .A(n74), .Y(n115) );
  INVX1 U81 ( .A(n80), .Y(n112) );
  INVX1 U82 ( .A(n75), .Y(n113) );
  INVX1 U83 ( .A(n79), .Y(n110) );
  INVX1 U84 ( .A(n88), .Y(n111) );
  INVX1 U85 ( .A(n89), .Y(n102) );
  INVX1 U86 ( .A(n78), .Y(n101) );
  INVX1 U87 ( .A(n84), .Y(n120) );
  INVX1 U88 ( .A(n71), .Y(n121) );
  INVX1 U89 ( .A(r_avg00[9]), .Y(n38) );
  INVX1 U90 ( .A(n35), .Y(dacyc_done) );
  INVX1 U91 ( .A(r_avg00[0]), .Y(n47) );
  INVX1 U92 ( .A(r_avg00[1]), .Y(n46) );
  INVX1 U93 ( .A(r_avg00[2]), .Y(n45) );
  INVX1 U94 ( .A(r_avg00[3]), .Y(n44) );
  INVX1 U95 ( .A(r_avg00[4]), .Y(n43) );
  INVX1 U96 ( .A(r_avg00[5]), .Y(n42) );
  INVX1 U97 ( .A(r_avg00[6]), .Y(n41) );
  INVX1 U98 ( .A(r_avg00[7]), .Y(n40) );
  INVX1 U99 ( .A(n65), .Y(sacyc_done) );
  INVX1 U100 ( .A(n70), .Y(n123) );
  INVX1 U101 ( .A(n85), .Y(n122) );
  INVX1 U102 ( .A(n23), .Y(n21) );
  INVX1 U103 ( .A(n23), .Y(n22) );
  INVX1 U104 ( .A(n86), .Y(n94) );
  AO21XL U105 ( .B(sar_nxt), .C(n23), .A(n8), .Y(updup) );
  MUX2X1 U106 ( .D0(n66), .D1(n67), .S(sarcyc[2]), .Y(N63) );
  AND2X1 U107 ( .A(n59), .B(n69), .Y(n66) );
  ENOX1 U108 ( .A(n11), .B(n88), .C(N88), .D(n11), .Y(rpt_v[6]) );
  OA21X1 U109 ( .B(sarcyc[1]), .C(sarcyc[0]), .A(n67), .Y(N62) );
  AND2X1 U110 ( .A(N42), .B(n49), .Y(N50) );
  AND2X1 U111 ( .A(N36), .B(n49), .Y(N44) );
  OAI22X1 U112 ( .A(n54), .B(n53), .C(n60), .D(n52), .Y(N64) );
  MUX2X1 U113 ( .D0(n52), .D1(n51), .S(sarcyc[2]), .Y(n54) );
  INVX1 U114 ( .A(sarcyc[3]), .Y(n52) );
  NAND21X1 U115 ( .B(sarcyc[3]), .A(n59), .Y(n51) );
  ENOX1 U116 ( .A(n124), .B(n91), .C(n124), .D(N91), .Y(rpt_v[9]) );
  ENOX1 U117 ( .A(n11), .B(n90), .C(N90), .D(n124), .Y(rpt_v[8]) );
  ENOX1 U118 ( .A(dac_v[0]), .B(n71), .C(N83), .D(n124), .Y(rpt_v[1]) );
  ENOX1 U119 ( .A(n124), .B(n72), .C(N84), .D(n124), .Y(rpt_v[2]) );
  ENOX1 U120 ( .A(n11), .B(n75), .C(N87), .D(n11), .Y(rpt_v[5]) );
  ENOX1 U121 ( .A(n124), .B(n73), .C(N85), .D(n11), .Y(rpt_v[3]) );
  ENOX1 U122 ( .A(n124), .B(n74), .C(N86), .D(n124), .Y(rpt_v[4]) );
  ENOX1 U123 ( .A(n11), .B(n89), .C(N89), .D(n11), .Y(rpt_v[7]) );
  ENOX1 U124 ( .A(n11), .B(n70), .C(N82), .D(n11), .Y(rpt_v[0]) );
  XNOR2XL U125 ( .A(dacnt[6]), .B(N23), .Y(n63) );
  XNOR2XL U126 ( .A(dacnt[3]), .B(N20), .Y(n62) );
  XOR2X1 U127 ( .A(dacnt[5]), .B(N23), .Y(n58) );
  NOR3XL U128 ( .A(n57), .B(n55), .C(n56), .Y(sampl_done) );
  NAND2X1 U129 ( .A(n58), .B(n92), .Y(n56) );
  NAND4X1 U130 ( .A(dacnt[1]), .B(n61), .C(n62), .D(n63), .Y(n55) );
  XOR2X1 U131 ( .A(N21), .B(dacnt[4]), .Y(n57) );
  AOI21X1 U132 ( .B(r_dac_t[0]), .C(r_dac_t[1]), .A(n107), .Y(N20) );
  OAI21X1 U133 ( .B(r_dac_t[0]), .C(n107), .A(n93), .Y(N21) );
  NOR2X1 U134 ( .A(r_dac_t[1]), .B(r_dac_t[0]), .Y(n107) );
  XNOR2XL U135 ( .A(dacnt[2]), .B(N19), .Y(n61) );
  NOR2X1 U136 ( .A(n107), .B(r_dac_t[1]), .Y(N19) );
  INVX1 U137 ( .A(dacnt[0]), .Y(n92) );
  NAND42X1 U138 ( .C(dacnt[1]), .D(dacnt[2]), .A(n86), .B(n87), .Y(n64) );
  NOR4XL U139 ( .A(dacnt[6]), .B(dacnt[5]), .C(dacnt[4]), .D(dacnt[3]), .Y(n87) );
  MUX2AXL U140 ( .D0(r_lt_lo[8]), .D1(n39), .S(n21), .Y(n77) );
  MUX2BXL U141 ( .D0(n45), .D1(r_lt_up[2]), .S(n22), .Y(n72) );
  MUX2BXL U142 ( .D0(n44), .D1(r_lt_up[3]), .S(n22), .Y(n73) );
  MUX2BXL U143 ( .D0(n43), .D1(r_lt_up[4]), .S(n22), .Y(n74) );
  MUX2BXL U144 ( .D0(n42), .D1(r_lt_up[5]), .S(n22), .Y(n75) );
  MUX2BXL U145 ( .D0(n41), .D1(r_lt_up[6]), .S(n22), .Y(n88) );
  MUX2BXL U146 ( .D0(n40), .D1(r_lt_up[7]), .S(n22), .Y(n89) );
  MUX2BXL U147 ( .D0(n39), .D1(r_lt_up[8]), .S(n22), .Y(n90) );
  MUX2BXL U148 ( .D0(n38), .D1(r_lt_up[9]), .S(n21), .Y(n91) );
  MUX2BXL U149 ( .D0(n47), .D1(r_lt_up[0]), .S(n22), .Y(n70) );
  MUX2BXL U150 ( .D0(n46), .D1(r_lt_up[1]), .S(n22), .Y(n71) );
  MUX2AXL U151 ( .D0(r_lt_lo[0]), .D1(n47), .S(n22), .Y(n85) );
  MUX2AXL U152 ( .D0(r_lt_lo[1]), .D1(n46), .S(n21), .Y(n84) );
  MUX2AXL U153 ( .D0(r_lt_lo[2]), .D1(n45), .S(n21), .Y(n83) );
  MUX2AXL U154 ( .D0(r_lt_lo[3]), .D1(n44), .S(n21), .Y(n82) );
  MUX2AXL U155 ( .D0(r_lt_lo[4]), .D1(n43), .S(n21), .Y(n81) );
  MUX2AXL U156 ( .D0(r_lt_lo[5]), .D1(n42), .S(n21), .Y(n80) );
  MUX2AXL U157 ( .D0(r_lt_lo[6]), .D1(n41), .S(n21), .Y(n79) );
  MUX2AXL U158 ( .D0(r_lt_lo[7]), .D1(n40), .S(n21), .Y(n78) );
  MUX2AXL U159 ( .D0(r_lt_lo[9]), .D1(n38), .S(n21), .Y(n76) );
  NAND32X1 U160 ( .B(n98), .C(n97), .A(n32), .Y(n65) );
  XNOR2XL U161 ( .A(sarcyc[2]), .B(r_sar10), .Y(n98) );
  XNOR2XL U162 ( .A(sarcyc[1]), .B(r_sar10), .Y(n97) );
  AND3X1 U163 ( .A(sarcyc[0]), .B(dacyc_done), .C(n31), .Y(n32) );
  NAND43X1 U164 ( .B(n104), .C(n103), .D(n105), .A(n30), .Y(n35) );
  XNOR2XL U165 ( .A(dacnt[3]), .B(n108), .Y(n104) );
  AND4X1 U166 ( .A(dacnt[1]), .B(dacnt[0]), .C(n29), .D(n28), .Y(n30) );
  XNOR2XL U167 ( .A(dacnt[2]), .B(n109), .Y(n103) );
  XNOR2XL U168 ( .A(r_sar10), .B(sarcyc[3]), .Y(n31) );
  XNOR2XL U169 ( .A(dacnt[4]), .B(n106), .Y(n105) );
  AOI22X1 U170 ( .A(n86), .B(N21), .C(r_dacyc), .D(n94), .Y(n106) );
  XOR2X1 U171 ( .A(dacnt[6]), .B(n19), .Y(n28) );
  OR2X1 U172 ( .A(n93), .B(n94), .Y(n19) );
  XOR2X1 U173 ( .A(dacnt[5]), .B(n20), .Y(n29) );
  OR2X1 U174 ( .A(N23), .B(n94), .Y(n20) );
  AOI22X1 U175 ( .A(N19), .B(n86), .C(r_dacyc), .D(n94), .Y(n109) );
  EORX1 U176 ( .A(N20), .B(n86), .C(r_dacyc), .D(n86), .Y(n108) );
  INVX1 U177 ( .A(sync_i), .Y(n23) );
  INVX1 U178 ( .A(n50), .Y(n59) );
  NAND21X1 U179 ( .B(n68), .A(sarcyc[1]), .Y(n50) );
  INVX1 U180 ( .A(sarcyc[0]), .Y(n68) );
endmodule


module dac2sar_a0_DW01_add_3 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n6, n7, n8, n9, n18, n19, n21, n23, n24, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n37, n39, n40, n45, n46, n49, n50, n51,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n68,
         n70, n71, n72, n73, n74, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125;

  XOR2X1 U22 ( .A(n31), .B(n3), .Y(SUM[7]) );
  OAI21X1 U27 ( .B(n29), .C(n37), .A(n30), .Y(n28) );
  OAI21X1 U66 ( .B(n56), .C(n60), .A(n57), .Y(n55) );
  XOR2X1 U71 ( .A(n61), .B(n8), .Y(SUM[2]) );
  OAI21X1 U72 ( .B(n61), .C(n59), .A(n60), .Y(n58) );
  XOR2X1 U77 ( .A(n9), .B(n65), .Y(SUM[1]) );
  NOR2X1 U88 ( .A(A[6]), .B(B[6]), .Y(n34) );
  NOR2XL U89 ( .A(A[7]), .B(B[7]), .Y(n29) );
  INVX1 U90 ( .A(n23), .Y(n21) );
  NAND2XL U91 ( .A(A[8]), .B(B[8]), .Y(n23) );
  NOR2X1 U92 ( .A(A[3]), .B(B[3]), .Y(n56) );
  NOR2X1 U93 ( .A(n34), .B(n29), .Y(n27) );
  NAND2X1 U94 ( .A(A[0]), .B(B[0]), .Y(n65) );
  NOR2X1 U95 ( .A(A[1]), .B(B[1]), .Y(n63) );
  AO21XL U96 ( .B(n24), .C(n116), .A(n119), .Y(SUM[10]) );
  OR2X1 U97 ( .A(A[9]), .B(B[9]), .Y(n114) );
  AND2X1 U98 ( .A(n39), .B(n27), .Y(n115) );
  AND2X1 U99 ( .A(n120), .B(n114), .Y(n116) );
  NAND2XL U100 ( .A(A[1]), .B(B[1]), .Y(n64) );
  AOI21XL U101 ( .B(n117), .C(n32), .A(n33), .Y(n31) );
  NAND2X1 U102 ( .A(n118), .B(n26), .Y(n24) );
  NAND2X1 U103 ( .A(A[3]), .B(B[3]), .Y(n57) );
  NAND2XL U104 ( .A(n120), .B(n23), .Y(n2) );
  XNOR2XL U105 ( .A(n2), .B(n24), .Y(SUM[8]) );
  OR2X1 U106 ( .A(A[8]), .B(B[8]), .Y(n120) );
  NAND2X1 U107 ( .A(n117), .B(n115), .Y(n118) );
  INVXL U108 ( .A(n53), .Y(n117) );
  AOI21X1 U109 ( .B(n27), .C(n40), .A(n28), .Y(n26) );
  AOI21XL U110 ( .B(n54), .C(n62), .A(n55), .Y(n53) );
  INVXL U111 ( .A(n51), .Y(n49) );
  NOR2XL U112 ( .A(A[5]), .B(B[5]), .Y(n45) );
  NOR2XL U113 ( .A(A[4]), .B(B[4]), .Y(n50) );
  NAND2XL U114 ( .A(A[5]), .B(B[5]), .Y(n46) );
  NAND2X1 U115 ( .A(n114), .B(n18), .Y(n1) );
  XOR2XL U116 ( .A(n123), .B(n124), .Y(SUM[6]) );
  XOR2XL U117 ( .A(n121), .B(n122), .Y(SUM[5]) );
  OAI21BXL U118 ( .C(n40), .B(n34), .A(n37), .Y(n33) );
  OAI21BBX1 U119 ( .A(n114), .B(n21), .C(n18), .Y(n119) );
  NOR2X1 U120 ( .A(n50), .B(n45), .Y(n39) );
  INVXL U121 ( .A(n56), .Y(n72) );
  INVXL U122 ( .A(n29), .Y(n68) );
  INVX1 U123 ( .A(n50), .Y(n71) );
  NOR21XL U124 ( .B(n39), .A(n34), .Y(n32) );
  NOR2X1 U125 ( .A(A[2]), .B(B[2]), .Y(n59) );
  NAND2XL U126 ( .A(A[9]), .B(B[9]), .Y(n18) );
  NAND2X1 U127 ( .A(A[6]), .B(B[6]), .Y(n37) );
  NAND2X1 U128 ( .A(A[4]), .B(B[4]), .Y(n51) );
  NAND2X1 U129 ( .A(A[2]), .B(B[2]), .Y(n60) );
  OR2XL U130 ( .A(A[6]), .B(B[6]), .Y(n125) );
  NAND2XL U131 ( .A(A[7]), .B(B[7]), .Y(n30) );
  NAND2XL U132 ( .A(n68), .B(n30), .Y(n3) );
  AO21XL U133 ( .B(n117), .C(n71), .A(n49), .Y(n121) );
  AND2XL U134 ( .A(n70), .B(n46), .Y(n122) );
  NAND2XL U135 ( .A(n74), .B(n64), .Y(n9) );
  AO21XL U136 ( .B(n117), .C(n39), .A(n40), .Y(n123) );
  AND2XL U137 ( .A(n125), .B(n37), .Y(n124) );
  NAND2XL U138 ( .A(n73), .B(n60), .Y(n8) );
  INVXL U139 ( .A(n59), .Y(n73) );
  XNOR2XL U140 ( .A(n6), .B(n117), .Y(SUM[4]) );
  XNOR2XL U141 ( .A(n7), .B(n58), .Y(SUM[3]) );
  NAND2XL U142 ( .A(n72), .B(n57), .Y(n7) );
  OAI21X1 U143 ( .B(n45), .C(n51), .A(n46), .Y(n40) );
  INVX1 U144 ( .A(n45), .Y(n70) );
  NAND2X1 U145 ( .A(n71), .B(n51), .Y(n6) );
  INVXL U146 ( .A(n62), .Y(n61) );
  NOR2XL U147 ( .A(n59), .B(n56), .Y(n54) );
  INVXL U148 ( .A(n63), .Y(n74) );
  OAI21X1 U149 ( .B(n63), .C(n65), .A(n64), .Y(n62) );
  XOR2X1 U150 ( .A(n19), .B(n1), .Y(SUM[9]) );
  AOI21X1 U151 ( .B(n24), .C(n120), .A(n21), .Y(n19) );
endmodule


module dac2sar_a0_DW01_inc_0 ( A, SUM );
  input [6:0] A;
  output [6:0] SUM;

  wire   [6:2] carry;

  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  XOR2X1 U1 ( .A(carry[6]), .B(A[6]), .Y(SUM[6]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module dac2sar_a0_DW01_add_2 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;

  wire   [9:1] carry;

  FAD1X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(SUM[10]), .SO(SUM[9])
         );
  FAD1X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .SO(SUM[8])
         );
  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  AND2X1 U1 ( .A(B[0]), .B(A[0]), .Y(carry[1]) );
endmodule


module dac2sar_a0_DW01_add_0 ( A, B, CI, SUM, CO );
  input [10:0] A;
  input [10:0] B;
  output [10:0] SUM;
  input CI;
  output CO;

  wire   [9:1] carry;

  FAD1X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(SUM[10]), .SO(SUM[9])
         );
  FAD1X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .SO(SUM[8])
         );
  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  AND2X1 U1 ( .A(B[0]), .B(A[0]), .Y(carry[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dac2sar_a0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dac2sar_a0_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_WIDTH10_0 ( clk, arstz, we, wdat, rdat );
  input [9:0] wdat;
  output [9:0] rdat;
  input clk, arstz, we;
  wire   net10209;

  SNPS_CLOCK_GATE_HIGH_glreg_WIDTH10_0 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10209), .TE(1'b0) );
  DFFRQX1 mem_reg_9_ ( .D(wdat[9]), .C(net10209), .XR(arstz), .Q(rdat[9]) );
  DFFRQX1 mem_reg_8_ ( .D(wdat[8]), .C(net10209), .XR(arstz), .Q(rdat[8]) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net10209), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net10209), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net10209), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net10209), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net10209), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net10209), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net10209), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net10209), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_WIDTH10_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_WIDTH10_1 ( clk, arstz, we, wdat, rdat );
  input [9:0] wdat;
  output [9:0] rdat;
  input clk, arstz, we;
  wire   net10227;

  SNPS_CLOCK_GATE_HIGH_glreg_WIDTH10_1 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10227), .TE(1'b0) );
  DFFRQX1 mem_reg_9_ ( .D(wdat[9]), .C(net10227), .XR(arstz), .Q(rdat[9]) );
  DFFRQX1 mem_reg_8_ ( .D(wdat[8]), .C(net10227), .XR(arstz), .Q(rdat[8]) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net10227), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net10227), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net10227), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net10227), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net10227), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net10227), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net10227), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net10227), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_WIDTH10_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_WIDTH10_2 ( clk, arstz, we, wdat, rdat );
  input [9:0] wdat;
  output [9:0] rdat;
  input clk, arstz, we;
  wire   net10245;

  SNPS_CLOCK_GATE_HIGH_glreg_WIDTH10_2 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10245), .TE(1'b0) );
  DFFRQXL mem_reg_7_ ( .D(wdat[7]), .C(net10245), .XR(arstz), .Q(rdat[7]) );
  DFFRQXL mem_reg_4_ ( .D(wdat[4]), .C(net10245), .XR(arstz), .Q(rdat[4]) );
  DFFRQXL mem_reg_3_ ( .D(wdat[3]), .C(net10245), .XR(arstz), .Q(rdat[3]) );
  DFFRQXL mem_reg_2_ ( .D(wdat[2]), .C(net10245), .XR(arstz), .Q(rdat[2]) );
  DFFRQXL mem_reg_1_ ( .D(wdat[1]), .C(net10245), .XR(arstz), .Q(rdat[1]) );
  DFFRQXL mem_reg_9_ ( .D(wdat[9]), .C(net10245), .XR(arstz), .Q(rdat[9]) );
  DFFRQXL mem_reg_8_ ( .D(wdat[8]), .C(net10245), .XR(arstz), .Q(rdat[8]) );
  DFFRQXL mem_reg_6_ ( .D(wdat[6]), .C(net10245), .XR(arstz), .Q(rdat[6]) );
  DFFRQXL mem_reg_5_ ( .D(wdat[5]), .C(net10245), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net10245), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_WIDTH10_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_00000012 ( clk, arstz, we, wdat, rdat );
  input [17:0] wdat;
  output [17:0] rdat;
  input clk, arstz, we;
  wire   net10263, n1, n2, n3;

  SNPS_CLOCK_GATE_HIGH_glreg_00000012 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10263), .TE(1'b0) );
  DFFRQX1 mem_reg_14_ ( .D(wdat[14]), .C(net10263), .XR(n1), .Q(rdat[14]) );
  DFFRQX1 mem_reg_13_ ( .D(wdat[13]), .C(net10263), .XR(n1), .Q(rdat[13]) );
  DFFRQX1 mem_reg_11_ ( .D(wdat[11]), .C(net10263), .XR(n1), .Q(rdat[11]) );
  DFFRQX1 mem_reg_9_ ( .D(wdat[9]), .C(net10263), .XR(n1), .Q(rdat[9]) );
  DFFRQX1 mem_reg_17_ ( .D(wdat[17]), .C(net10263), .XR(n1), .Q(rdat[17]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net10263), .XR(n2), .Q(rdat[0]) );
  DFFRQX1 mem_reg_12_ ( .D(wdat[12]), .C(net10263), .XR(n1), .Q(rdat[12]) );
  DFFRQX1 mem_reg_10_ ( .D(wdat[10]), .C(net10263), .XR(n1), .Q(rdat[10]) );
  DFFRQX1 mem_reg_8_ ( .D(wdat[8]), .C(net10263), .XR(n1), .Q(rdat[8]) );
  DFFRQX1 mem_reg_16_ ( .D(wdat[16]), .C(net10263), .XR(n1), .Q(rdat[16]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net10263), .XR(n2), .Q(rdat[5]) );
  DFFRQX1 mem_reg_15_ ( .D(wdat[15]), .C(net10263), .XR(n1), .Q(rdat[15]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net10263), .XR(n2), .Q(rdat[6]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net10263), .XR(n2), .Q(rdat[4]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net10263), .XR(n2), .Q(rdat[2]) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net10263), .XR(n2), .Q(rdat[7]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net10263), .XR(n2), .Q(rdat[3]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net10263), .XR(n2), .Q(rdat[1]) );
  INVX1 U2 ( .A(n3), .Y(n1) );
  INVX1 U3 ( .A(n3), .Y(n2) );
  INVX1 U4 ( .A(arstz), .Y(n3) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_00000012 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module updphy_FF_DEPTH_NUM34_FF_DEPTH_NBT6 ( i_cc, i_cc_49, i_sqlch, r_sqlch, 
        r_adprx_en, r_adp2nd, r_exist1st, r_ordrs4, r_fifopsh, r_fifopop, 
        r_fiforst, r_unlock, r_first, r_last, r_set_cpmsgid, r_rdy, r_wdat, 
        r_rdat, r_txnumk, r_txendk, r_txshrt, r_auto_discard, r_txauto, 
        r_rxords_ena, r_spec, r_dat_spec, r_auto_gdcrc, r_rxdb_opt, r_pshords, 
        r_dat_portrole, r_dat_datarole, r_discard, pid_goidle, pid_gobusy, 
        pff_ack, pff_rdat, pff_rxpart, prx_rcvinf, pff_obsd, pff_ptr, 
        pff_empty, pff_full, ptx_ack, ptx_cc, ptx_oe, prx_setsta, prx_rst, 
        prl_c0set, prl_cany0, prl_cany0r, prl_cany0w, prl_discard, 
        prl_GCTxDone, prl_cany0adr, prl_cpmsgid, prx_fifowdat, ptx_fsm, 
        prl_fsm, prx_fsm, prx_adpn, dbgpo, clk, srstz );
  input [1:0] r_sqlch;
  input [7:0] r_wdat;
  input [7:0] r_rdat;
  input [4:0] r_txnumk;
  input [6:0] r_txauto;
  input [6:0] r_rxords_ena;
  input [1:0] r_spec;
  input [1:0] r_dat_spec;
  input [1:0] r_auto_gdcrc;
  input [1:0] r_rxdb_opt;
  output [1:0] pff_ack;
  output [7:0] pff_rdat;
  output [15:0] pff_rxpart;
  output [4:0] prx_rcvinf;
  output [5:0] pff_ptr;
  output [6:0] prx_setsta;
  output [1:0] prx_rst;
  output [7:0] prl_cany0adr;
  output [2:0] prl_cpmsgid;
  output [7:0] prx_fifowdat;
  output [2:0] ptx_fsm;
  output [3:0] prl_fsm;
  output [3:0] prx_fsm;
  output [5:0] prx_adpn;
  output [31:0] dbgpo;
  input i_cc, i_cc_49, i_sqlch, r_adprx_en, r_adp2nd, r_exist1st, r_ordrs4,
         r_fifopsh, r_fifopop, r_fiforst, r_unlock, r_first, r_last,
         r_set_cpmsgid, r_rdy, r_txendk, r_txshrt, r_auto_discard, r_pshords,
         r_dat_portrole, r_dat_datarole, r_discard, clk, srstz;
  output pid_goidle, pid_gobusy, pff_obsd, pff_empty, pff_full, ptx_ack,
         ptx_cc, ptx_oe, prl_c0set, prl_cany0, prl_cany0r, prl_cany0w,
         prl_discard, prl_GCTxDone;
  wire   n56, rx_pshords, auto_rx_gdcrc, prx_trans, prx_fiforst, pcc_rxgood,
         prx_crcstart, prx_crcshfi4, prx_eoprcvd, x_trans, ptx_goidle,
         c0_txendk, mux_one, ptx_crcstart, ptx_crcshfi4, ptx_crcshfo4,
         crcstart, crcshfi4, crcshfo4, prl_idle, lockena, fifosrstz,
         fifopop_pff, fifopsh_pff, pff_txreq, pff_one, obsd, prl_last,
         prl_txreq, fifopop_prl, fifopsh_prl, prx_gdmsgrcvd, N25, N26, N27,
         N28, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41,
         N42, N43, d_sqlch, net10281, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n3, n5, n6, n21, n22, n23, n24, n25, n26,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2,
         SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4;
  wire   [1:0] prx_cccnt;
  wire   [3:0] prx_crcsidat;
  wire   [4:0] c0_txnumk;
  wire   [6:0] c0_txauto;
  wire   [7:0] mux_rdat;
  wire   [3:0] ptx_crcsidat;
  wire   [3:0] crc32_3_0;
  wire   [3:0] crcsidat;
  wire   [55:0] pff_dat_7_1;
  wire   [47:16] pff_c0dat;
  wire   [7:0] prl_rdat;
  wire   [4:0] prl_txauto;
  wire   [1:0] d_cc;
  wire   [8:0] cclow_cnt;

  phyrx_a0 u0_phyrx ( .i_cc(i_cc), .ptx_txact(n5), .r_adprx_en(r_adprx_en), 
        .r_adp2nd(r_adp2nd), .r_exist1st(r_exist1st), .r_ordrs4(r_ordrs4), 
        .r_rxdb_opt(r_rxdb_opt), .r_ords_ena(r_rxords_ena), .r_pshords(
        rx_pshords), .r_rgdcrc(auto_rx_gdcrc), .prx_cccnt(prx_cccnt), 
        .prx_rst(prx_rst), .prx_setsta({prx_setsta[6:1], 
        SYNOPSYS_UNCONNECTED_1}), .prx_idle(), .prx_d_cc(prx_rcvinf[3]), 
        .prx_bmc(dbgpo[18]), .prx_trans(prx_trans), .prx_fiforst(prx_fiforst), 
        .prx_fifopsh(dbgpo[29]), .prx_fifowdat(prx_fifowdat), .pff_txreq(n6), 
        .pid_gobusy(pid_gobusy), .pid_goidle(pid_goidle), .pid_ccidle(
        prx_rcvinf[4]), .pcc_rxgood(pcc_rxgood), .prx_crcstart(prx_crcstart), 
        .prx_crcshfi4(prx_crcshfi4), .prx_crcsidat(prx_crcsidat), .prx_rxcode(
        dbgpo[28:24]), .prx_adpn(prx_adpn), .prx_rcvdords(prx_rcvinf[2:0]), 
        .prx_eoprcvd(prx_eoprcvd), .prx_fsm(prx_fsm), .clk(clk), .srstz(n25)
         );
  phyidd_a0 u0_phyidd ( .i_trans(x_trans), .i_goidle(ptx_goidle), .o_ccidle(
        prx_rcvinf[4]), .o_goidle(pid_goidle), .o_gobusy(pid_gobusy), .clk(clk), .srstz(n24) );
  phytx_a0 u0_phytx ( .r_txnumk(c0_txnumk), .r_txendk(c0_txendk), .r_txshrt(
        r_txshrt), .r_txauto(c0_txauto), .prx_cccnt(prx_cccnt), .ptx_txact(n56), .ptx_cc(ptx_cc), .ptx_goidle(ptx_goidle), .ptx_fifopop(dbgpo[30]), 
        .ptx_pspyld(), .i_rdat(mux_rdat), .i_txreq(n6), .i_one(mux_one), 
        .ptx_crcstart(ptx_crcstart), .ptx_crcshfi4(ptx_crcshfi4), 
        .ptx_crcshfo4(ptx_crcshfo4), .ptx_crcsidat(ptx_crcsidat), .ptx_fsm(
        ptx_fsm), .pcc_crc30(crc32_3_0), .clk(clk), .srstz(srstz) );
  phycrc_a0 u0_phycrc ( .crc32_3_0(crc32_3_0), .rx_good(pcc_rxgood), 
        .i_shfidat(crcsidat), .i_start(crcstart), .i_shfi4(crcshfi4), 
        .i_shfo4(crcshfo4), .clk(clk) );
  phyff_DEPTH_NUM34_DEPTH_NBT6 u0_phyff ( .r_psh(r_fifopsh), .r_pop(r_fifopop), 
        .prx_psh(fifopsh_pff), .ptx_pop(fifopop_pff), .r_last(r_last), 
        .r_unlock(r_unlock), .i_lockena(lockena), .r_fiforst(r_fiforst), 
        .i_ccidle(prx_rcvinf[4]), .r_wdat(r_wdat), .prx_wdat(prx_fifowdat), 
        .txreq(pff_txreq), .ffack(pff_ack), .rdat0(pff_rdat), .full(pff_full), 
        .empty(pff_empty), .one(pff_one), .half(), .obsd(obsd), .dat_7_1(
        pff_dat_7_1), .ptr(pff_ptr), .fifowdat(dbgpo[7:0]), .fifopsh(dbgpo[16]), .clk(clk), .srstz(fifosrstz) );
  updprl_a0 u0_updprl ( .r_spec(r_spec), .r_dat_spec(r_dat_spec), 
        .r_auto_txgdcrc(r_auto_gdcrc[0]), .r_dat_portrole(r_dat_portrole), 
        .r_dat_datarole(r_dat_datarole), .r_auto_discard(r_auto_discard), 
        .r_set_cpmsgid(r_set_cpmsgid), .r_dat_cpmsgid(r_wdat[2:0]), .r_rdat(
        r_rdat), .r_rdy(r_rdy), .pid_ccidle(prx_rcvinf[4]), .r_discard(
        r_discard), .ptx_ack(ptx_goidle), .ptx_txact(n5), .ptx_fifopop(
        fifopop_prl), .prx_fifopsh(fifopsh_prl), .prx_gdmsgrcvd(prx_gdmsgrcvd), 
        .prx_eoprcvd(prx_eoprcvd), .prx_rcvdords(prx_rcvinf[2:0]), 
        .prx_fifowdat(prx_fifowdat), .pff_c0dat({pff_c0dat, pff_rxpart}), 
        .prl_rdat(prl_rdat), .prl_txauto({SYNOPSYS_UNCONNECTED_2, 
        SYNOPSYS_UNCONNECTED_3, prl_txauto[4], SYNOPSYS_UNCONNECTED_4, 
        prl_txauto[2:0]}), .prl_last(prl_last), .prl_txreq(prl_txreq), 
        .prl_c0set(prl_c0set), .prl_cany0(prl_cany0), .prl_cany0r(prl_cany0r), 
        .prl_cany0w(prl_cany0w), .prl_idle(prl_idle), .prl_discard(prl_discard), .prl_GCTxDone(prl_GCTxDone), .prl_fsm(prl_fsm), .prl_cpmsgid(prl_cpmsgid), 
        .prl_cany0adr(prl_cany0adr), .clk(clk), .srstz(n24) );
  dbnc_WIDTH3 u0_sqlch_db ( .o_dbc(d_sqlch), .o_chg(), .i_org(i_sqlch), .clk(
        clk), .rstz(n24) );
  SNPS_CLOCK_GATE_HIGH_updphy_FF_DEPTH_NUM34_FF_DEPTH_NBT6 clk_gate_cclow_cnt_reg ( 
        .CLK(clk), .EN(N34), .ENCLK(net10281), .TE(1'b0) );
  DFFSQX1 d_cc_reg_1_ ( .D(d_cc[0]), .C(clk), .XS(n25), .Q(d_cc[1]) );
  DFFSQX1 d_cc_reg_0_ ( .D(i_cc_49), .C(clk), .XS(n25), .Q(d_cc[0]) );
  DFFQX1 cclow_cnt_reg_2_ ( .D(N37), .C(net10281), .Q(cclow_cnt[2]) );
  DFFQX1 cclow_cnt_reg_3_ ( .D(N38), .C(net10281), .Q(cclow_cnt[3]) );
  DFFQX1 cclow_cnt_reg_4_ ( .D(N39), .C(net10281), .Q(cclow_cnt[4]) );
  DFFQX1 cclow_cnt_reg_5_ ( .D(N40), .C(net10281), .Q(cclow_cnt[5]) );
  DFFQX1 cclow_cnt_reg_6_ ( .D(N41), .C(net10281), .Q(cclow_cnt[6]) );
  DFFQX1 cclow_cnt_reg_8_ ( .D(N43), .C(net10281), .Q(cclow_cnt[8]) );
  DFFQX1 cclow_cnt_reg_7_ ( .D(N42), .C(net10281), .Q(cclow_cnt[7]) );
  DFFQX1 cclow_cnt_reg_1_ ( .D(N36), .C(net10281), .Q(cclow_cnt[1]) );
  DFFQX1 cclow_cnt_reg_0_ ( .D(N35), .C(net10281), .Q(cclow_cnt[0]) );
  INVX1 U3 ( .A(1'b1), .Y(dbgpo[31]) );
  MUX2X1 U5 ( .D0(prl_rdat[6]), .D1(pff_rdat[6]), .S(n22), .Y(mux_rdat[6]) );
  MUX2X1 U6 ( .D0(prl_rdat[3]), .D1(pff_rdat[3]), .S(n21), .Y(mux_rdat[3]) );
  MUX2X1 U7 ( .D0(prl_rdat[7]), .D1(pff_rdat[7]), .S(n22), .Y(mux_rdat[7]) );
  MUX2X1 U8 ( .D0(prl_rdat[4]), .D1(pff_rdat[4]), .S(n21), .Y(mux_rdat[4]) );
  AND2X1 U9 ( .A(n44), .B(n22), .Y(rx_pshords) );
  AND2X1 U10 ( .A(dbgpo[30]), .B(n23), .Y(fifopop_prl) );
  INVX1 U11 ( .A(n56), .Y(n3) );
  INVX1 U12 ( .A(n3), .Y(ptx_oe) );
  INVX1 U13 ( .A(n3), .Y(n5) );
  BUFX3 U14 ( .A(prx_fsm[3]), .Y(dbgpo[23]) );
  BUFX3 U15 ( .A(prx_rcvinf[4]), .Y(dbgpo[19]) );
  BUFX3 U16 ( .A(prx_fsm[0]), .Y(dbgpo[20]) );
  BUFX3 U17 ( .A(prx_fsm[2]), .Y(dbgpo[22]) );
  BUFX3 U18 ( .A(prx_fsm[1]), .Y(dbgpo[21]) );
  BUFX3 U19 ( .A(pff_rdat[5]), .Y(dbgpo[13]) );
  BUFX3 U20 ( .A(pff_rdat[2]), .Y(dbgpo[10]) );
  BUFX3 U21 ( .A(pff_rdat[3]), .Y(dbgpo[11]) );
  BUFX3 U22 ( .A(pff_rdat[4]), .Y(dbgpo[12]) );
  BUFX3 U23 ( .A(pff_rdat[6]), .Y(dbgpo[14]) );
  BUFX3 U24 ( .A(pff_rdat[7]), .Y(dbgpo[15]) );
  BUFX3 U25 ( .A(pff_rdat[0]), .Y(dbgpo[8]) );
  BUFX3 U26 ( .A(pff_rdat[1]), .Y(dbgpo[9]) );
  AND2X1 U27 ( .A(r_txnumk[2]), .B(n22), .Y(c0_txnumk[2]) );
  AND2X1 U28 ( .A(r_txnumk[1]), .B(n21), .Y(c0_txnumk[1]) );
  AND2XL U29 ( .A(r_txnumk[3]), .B(n22), .Y(c0_txnumk[3]) );
  AND2XL U30 ( .A(dbgpo[30]), .B(n22), .Y(fifopop_pff) );
  MUX2XL U31 ( .D0(prl_last), .D1(pff_one), .S(n21), .Y(mux_one) );
  MUX2XL U32 ( .D0(prl_txreq), .D1(pff_txreq), .S(prl_idle), .Y(n6) );
  AND2XL U33 ( .A(dbgpo[29]), .B(n22), .Y(fifopsh_pff) );
  MUX2XL U34 ( .D0(pff_rdat[6]), .D1(pff_dat_7_1[14]), .S(n44), .Y(
        pff_rxpart[6]) );
  MUX2XL U35 ( .D0(pff_rdat[7]), .D1(pff_dat_7_1[15]), .S(n44), .Y(
        pff_rxpart[7]) );
  MUX2XL U36 ( .D0(pff_rdat[0]), .D1(pff_dat_7_1[8]), .S(n40), .Y(
        pff_rxpart[0]) );
  MUX2XL U37 ( .D0(pff_rdat[1]), .D1(pff_dat_7_1[9]), .S(n41), .Y(
        pff_rxpart[1]) );
  MUX2XL U38 ( .D0(pff_rdat[2]), .D1(pff_dat_7_1[10]), .S(n42), .Y(
        pff_rxpart[2]) );
  MUX2XL U39 ( .D0(pff_rdat[3]), .D1(pff_dat_7_1[11]), .S(n43), .Y(
        pff_rxpart[3]) );
  MUX2XL U40 ( .D0(pff_rdat[4]), .D1(pff_dat_7_1[12]), .S(n44), .Y(
        pff_rxpart[4]) );
  INVX1 U41 ( .A(n23), .Y(n21) );
  INVX1 U42 ( .A(n23), .Y(n22) );
  INVX1 U43 ( .A(prl_idle), .Y(n23) );
  AND2X1 U44 ( .A(prx_setsta[3]), .B(n28), .Y(prx_gdmsgrcvd) );
  NOR2X1 U45 ( .A(prx_fiforst), .B(n26), .Y(fifosrstz) );
  NOR21XL U46 ( .B(ptx_crcshfo4), .A(n3), .Y(crcshfo4) );
  INVX1 U47 ( .A(n26), .Y(n25) );
  AND2X2 U48 ( .A(dbgpo[29]), .B(n23), .Y(fifopsh_prl) );
  INVX1 U49 ( .A(n45), .Y(n44) );
  AO22X1 U50 ( .A(ptx_crcstart), .B(n5), .C(prx_crcstart), .D(n3), .Y(crcstart) );
  AO22X1 U51 ( .A(ptx_crcshfi4), .B(ptx_oe), .C(prx_crcshfi4), .D(n3), .Y(
        crcshfi4) );
  NOR21XL U52 ( .B(obsd), .A(prx_setsta[6]), .Y(pff_obsd) );
  NAND42X1 U53 ( .C(pff_rxpart[1]), .D(pff_rxpart[15]), .A(n29), .B(n30), .Y(
        n28) );
  NOR3XL U54 ( .A(pff_rxpart[2]), .B(pff_rxpart[4]), .C(pff_rxpart[3]), .Y(n29) );
  NOR41XL U55 ( .D(pff_rxpart[0]), .A(pff_rxpart[14]), .B(pff_rxpart[13]), .C(
        pff_rxpart[12]), .Y(n30) );
  INVX1 U56 ( .A(n45), .Y(n40) );
  INVX1 U57 ( .A(n45), .Y(n41) );
  INVX1 U58 ( .A(n45), .Y(n43) );
  INVX1 U59 ( .A(n45), .Y(n42) );
  INVX1 U60 ( .A(srstz), .Y(n26) );
  NAND21X1 U61 ( .B(n36), .A(n35), .Y(n33) );
  INVX1 U62 ( .A(n34), .Y(n54) );
  NAND3X1 U63 ( .A(n34), .B(n33), .C(n35), .Y(N34) );
  INVX1 U64 ( .A(n26), .Y(n24) );
  MUX2X1 U65 ( .D0(prl_rdat[5]), .D1(pff_rdat[5]), .S(n21), .Y(mux_rdat[5]) );
  MUX2X2 U66 ( .D0(prl_rdat[2]), .D1(pff_rdat[2]), .S(prl_idle), .Y(
        mux_rdat[2]) );
  MUX2XL U67 ( .D0(prl_rdat[1]), .D1(pff_rdat[1]), .S(n21), .Y(mux_rdat[1]) );
  AND2XL U68 ( .A(r_txnumk[0]), .B(n21), .Y(c0_txnumk[0]) );
  AND2XL U69 ( .A(r_txendk), .B(n21), .Y(c0_txendk) );
  AND2XL U70 ( .A(r_txnumk[4]), .B(n22), .Y(c0_txnumk[4]) );
  MUX2XL U71 ( .D0(prl_rdat[0]), .D1(pff_rdat[0]), .S(n21), .Y(mux_rdat[0]) );
  AND2XL U72 ( .A(r_txauto[6]), .B(n21), .Y(c0_txauto[6]) );
  INVX1 U73 ( .A(r_pshords), .Y(n45) );
  AOI21AXL U74 ( .B(n5), .C(n22), .A(r_first), .Y(lockena) );
  NAND21XL U75 ( .B(r_txauto[5]), .A(prl_idle), .Y(c0_txauto[5]) );
  AO22X1 U76 ( .A(ptx_crcsidat[1]), .B(n5), .C(prx_crcsidat[1]), .D(n3), .Y(
        crcsidat[1]) );
  AO22XL U77 ( .A(ptx_crcsidat[3]), .B(n5), .C(prx_crcsidat[3]), .D(n3), .Y(
        crcsidat[3]) );
  MUX2X1 U78 ( .D0(pff_dat_7_1[8]), .D1(pff_dat_7_1[24]), .S(n40), .Y(
        pff_c0dat[16]) );
  MUX2X1 U79 ( .D0(pff_dat_7_1[10]), .D1(pff_dat_7_1[26]), .S(n40), .Y(
        pff_c0dat[18]) );
  MUX2X1 U80 ( .D0(pff_dat_7_1[16]), .D1(pff_dat_7_1[32]), .S(n41), .Y(
        pff_c0dat[24]) );
  MUX2X1 U81 ( .D0(pff_dat_7_1[13]), .D1(pff_dat_7_1[29]), .S(n41), .Y(
        pff_c0dat[21]) );
  MUX2X1 U82 ( .D0(pff_rdat[5]), .D1(pff_dat_7_1[13]), .S(n44), .Y(
        pff_rxpart[5]) );
  MUX2X1 U83 ( .D0(pff_dat_7_1[0]), .D1(pff_dat_7_1[16]), .S(n44), .Y(
        pff_rxpart[8]) );
  MUX2X1 U84 ( .D0(pff_dat_7_1[4]), .D1(pff_dat_7_1[20]), .S(n40), .Y(
        pff_rxpart[12]) );
  MUX2X1 U85 ( .D0(pff_dat_7_1[5]), .D1(pff_dat_7_1[21]), .S(n40), .Y(
        pff_rxpart[13]) );
  MUX2X1 U86 ( .D0(pff_dat_7_1[6]), .D1(pff_dat_7_1[22]), .S(n40), .Y(
        pff_rxpart[14]) );
  MUX2X1 U87 ( .D0(pff_dat_7_1[7]), .D1(pff_dat_7_1[23]), .S(n40), .Y(
        pff_rxpart[15]) );
  NOR21XL U88 ( .B(r_auto_gdcrc[1]), .A(n28), .Y(auto_rx_gdcrc) );
  MUX2X1 U89 ( .D0(pff_dat_7_1[39]), .D1(pff_dat_7_1[55]), .S(n44), .Y(
        pff_c0dat[47]) );
  MUX2X1 U90 ( .D0(pff_dat_7_1[37]), .D1(pff_dat_7_1[53]), .S(n43), .Y(
        pff_c0dat[45]) );
  MUX2X1 U91 ( .D0(pff_dat_7_1[11]), .D1(pff_dat_7_1[27]), .S(n41), .Y(
        pff_c0dat[19]) );
  MUX2X1 U92 ( .D0(pff_dat_7_1[34]), .D1(pff_dat_7_1[50]), .S(n43), .Y(
        pff_c0dat[42]) );
  MUX2X1 U93 ( .D0(pff_dat_7_1[25]), .D1(pff_dat_7_1[41]), .S(n42), .Y(
        pff_c0dat[33]) );
  MUX2X1 U94 ( .D0(pff_dat_7_1[22]), .D1(pff_dat_7_1[38]), .S(n42), .Y(
        pff_c0dat[30]) );
  MUX2X1 U95 ( .D0(pff_dat_7_1[32]), .D1(pff_dat_7_1[48]), .S(n43), .Y(
        pff_c0dat[40]) );
  MUX2X1 U96 ( .D0(pff_dat_7_1[29]), .D1(pff_dat_7_1[45]), .S(n43), .Y(
        pff_c0dat[37]) );
  MUX2X1 U97 ( .D0(pff_dat_7_1[27]), .D1(pff_dat_7_1[43]), .S(n42), .Y(
        pff_c0dat[35]) );
  MUX2X1 U98 ( .D0(pff_dat_7_1[38]), .D1(pff_dat_7_1[54]), .S(n44), .Y(
        pff_c0dat[46]) );
  MUX2X1 U99 ( .D0(pff_dat_7_1[28]), .D1(pff_dat_7_1[44]), .S(n42), .Y(
        pff_c0dat[36]) );
  MUX2X1 U100 ( .D0(pff_dat_7_1[14]), .D1(pff_dat_7_1[30]), .S(n41), .Y(
        pff_c0dat[22]) );
  MUX2X1 U101 ( .D0(pff_dat_7_1[26]), .D1(pff_dat_7_1[42]), .S(n42), .Y(
        pff_c0dat[34]) );
  MUX2X1 U102 ( .D0(pff_dat_7_1[12]), .D1(pff_dat_7_1[28]), .S(n41), .Y(
        pff_c0dat[20]) );
  MUX2X1 U103 ( .D0(pff_dat_7_1[9]), .D1(pff_dat_7_1[25]), .S(n40), .Y(
        pff_c0dat[17]) );
  MUX2X1 U104 ( .D0(pff_dat_7_1[35]), .D1(pff_dat_7_1[51]), .S(n43), .Y(
        pff_c0dat[43]) );
  MUX2X1 U105 ( .D0(pff_dat_7_1[23]), .D1(pff_dat_7_1[39]), .S(n42), .Y(
        pff_c0dat[31]) );
  MUX2X1 U106 ( .D0(pff_dat_7_1[21]), .D1(pff_dat_7_1[37]), .S(n42), .Y(
        pff_c0dat[29]) );
  MUX2X1 U107 ( .D0(pff_dat_7_1[36]), .D1(pff_dat_7_1[52]), .S(n43), .Y(
        pff_c0dat[44]) );
  MUX2X1 U108 ( .D0(pff_dat_7_1[24]), .D1(pff_dat_7_1[40]), .S(n42), .Y(
        pff_c0dat[32]) );
  MUX2X1 U109 ( .D0(pff_dat_7_1[33]), .D1(pff_dat_7_1[49]), .S(n43), .Y(
        pff_c0dat[41]) );
  MUX2X1 U110 ( .D0(pff_dat_7_1[31]), .D1(pff_dat_7_1[47]), .S(n43), .Y(
        pff_c0dat[39]) );
  MUX2X1 U111 ( .D0(pff_dat_7_1[30]), .D1(pff_dat_7_1[46]), .S(n43), .Y(
        pff_c0dat[38]) );
  MUX2X1 U112 ( .D0(pff_dat_7_1[18]), .D1(pff_dat_7_1[34]), .S(n41), .Y(
        pff_c0dat[26]) );
  MUX2X1 U113 ( .D0(pff_dat_7_1[17]), .D1(pff_dat_7_1[33]), .S(n41), .Y(
        pff_c0dat[25]) );
  MUX2X1 U114 ( .D0(pff_dat_7_1[15]), .D1(pff_dat_7_1[31]), .S(n41), .Y(
        pff_c0dat[23]) );
  MUX2X1 U115 ( .D0(pff_dat_7_1[20]), .D1(pff_dat_7_1[36]), .S(n42), .Y(
        pff_c0dat[28]) );
  MUX2X1 U116 ( .D0(pff_dat_7_1[19]), .D1(pff_dat_7_1[35]), .S(n41), .Y(
        pff_c0dat[27]) );
  MUX2XL U117 ( .D0(prl_txauto[0]), .D1(r_txauto[0]), .S(prl_idle), .Y(
        c0_txauto[0]) );
  MUX2XL U118 ( .D0(prl_txauto[2]), .D1(r_txauto[2]), .S(prl_idle), .Y(
        c0_txauto[2]) );
  MUX2XL U119 ( .D0(prl_txauto[1]), .D1(r_txauto[1]), .S(prl_idle), .Y(
        c0_txauto[1]) );
  MUX2XL U120 ( .D0(prl_txauto[4]), .D1(r_txauto[4]), .S(prl_idle), .Y(
        c0_txauto[4]) );
  NOR21XL U121 ( .B(ptx_goidle), .A(prl_cany0), .Y(ptx_ack) );
  AOI31X1 U122 ( .A(d_sqlch), .B(n27), .C(r_sqlch[0]), .D(n53), .Y(x_trans) );
  INVX1 U123 ( .A(prx_trans), .Y(n53) );
  OAI21X1 U124 ( .B(prx_fsm[3]), .C(n5), .A(r_sqlch[1]), .Y(n27) );
  NAND21XL U125 ( .B(r_txauto[3]), .A(prl_idle), .Y(c0_txauto[3]) );
  OAI21BBX1 U126 ( .A(N33), .B(n54), .C(n33), .Y(N43) );
  NOR4XL U127 ( .A(n31), .B(n32), .C(cclow_cnt[5]), .D(cclow_cnt[4]), .Y(
        prx_setsta[0]) );
  OR3XL U128 ( .A(cclow_cnt[7]), .B(cclow_cnt[8]), .C(cclow_cnt[6]), .Y(n32)
         );
  NAND43X1 U129 ( .B(cclow_cnt[1]), .C(cclow_cnt[3]), .D(cclow_cnt[2]), .A(
        cclow_cnt[0]), .Y(n31) );
  AND2X1 U130 ( .A(N32), .B(n54), .Y(N42) );
  OAI21BBX1 U131 ( .A(N31), .B(n54), .C(n33), .Y(N41) );
  AOI21BBXL U132 ( .B(d_cc[1]), .C(n55), .A(n26), .Y(n35) );
  OAI211X1 U133 ( .C(n37), .D(n38), .A(n36), .B(n35), .Y(n34) );
  OR4X1 U134 ( .A(cclow_cnt[0]), .B(cclow_cnt[1]), .C(cclow_cnt[2]), .D(
        cclow_cnt[3]), .Y(n38) );
  NAND43X1 U135 ( .B(cclow_cnt[4]), .C(cclow_cnt[5]), .D(cclow_cnt[6]), .A(n39), .Y(n37) );
  NOR2X1 U136 ( .A(cclow_cnt[8]), .B(cclow_cnt[7]), .Y(n39) );
  AND2X1 U137 ( .A(N25), .B(n54), .Y(N35) );
  AND2X1 U138 ( .A(N28), .B(n54), .Y(N38) );
  AND2X1 U139 ( .A(N27), .B(n54), .Y(N37) );
  OAI21BBX1 U140 ( .A(N30), .B(n54), .C(n33), .Y(N40) );
  OAI21BBX1 U141 ( .A(N29), .B(n54), .C(n33), .Y(N39) );
  OAI21BBX1 U142 ( .A(N26), .B(n54), .C(n33), .Y(N36) );
  MUX2X1 U143 ( .D0(pff_dat_7_1[1]), .D1(pff_dat_7_1[17]), .S(n44), .Y(
        pff_rxpart[9]) );
  MUX2X1 U144 ( .D0(pff_dat_7_1[2]), .D1(pff_dat_7_1[18]), .S(n40), .Y(
        pff_rxpart[10]) );
  MUX2X1 U145 ( .D0(pff_dat_7_1[3]), .D1(pff_dat_7_1[19]), .S(n40), .Y(
        pff_rxpart[11]) );
  NAND2X1 U146 ( .A(d_cc[1]), .B(n55), .Y(n36) );
  INVX1 U147 ( .A(d_cc[0]), .Y(n55) );
  BUFX3 U148 ( .A(prx_rcvinf[3]), .Y(dbgpo[17]) );
  AO22XL U149 ( .A(ptx_crcsidat[2]), .B(n5), .C(prx_crcsidat[2]), .D(n3), .Y(
        crcsidat[2]) );
  AO22XL U150 ( .A(ptx_crcsidat[0]), .B(n5), .C(prx_crcsidat[0]), .D(n3), .Y(
        crcsidat[0]) );
  INVX1 U151 ( .A(cclow_cnt[0]), .Y(N25) );
  OR2X1 U152 ( .A(cclow_cnt[1]), .B(cclow_cnt[0]), .Y(n46) );
  OAI21BBX1 U153 ( .A(cclow_cnt[0]), .B(cclow_cnt[1]), .C(n46), .Y(N26) );
  OR2X1 U154 ( .A(n46), .B(cclow_cnt[2]), .Y(n47) );
  OAI21BBX1 U155 ( .A(n46), .B(cclow_cnt[2]), .C(n47), .Y(N27) );
  OR2X1 U156 ( .A(n47), .B(cclow_cnt[3]), .Y(n48) );
  OAI21BBX1 U157 ( .A(n47), .B(cclow_cnt[3]), .C(n48), .Y(N28) );
  OR2X1 U158 ( .A(n48), .B(cclow_cnt[4]), .Y(n49) );
  OAI21BBX1 U159 ( .A(n48), .B(cclow_cnt[4]), .C(n49), .Y(N29) );
  OR2X1 U160 ( .A(n49), .B(cclow_cnt[5]), .Y(n50) );
  OAI21BBX1 U161 ( .A(n49), .B(cclow_cnt[5]), .C(n50), .Y(N30) );
  OR2X1 U162 ( .A(n50), .B(cclow_cnt[6]), .Y(n51) );
  OAI21BBX1 U163 ( .A(n50), .B(cclow_cnt[6]), .C(n51), .Y(N31) );
  XNOR2XL U164 ( .A(n51), .B(cclow_cnt[7]), .Y(N32) );
  OR2X1 U165 ( .A(cclow_cnt[7]), .B(n51), .Y(n52) );
  XNOR2XL U166 ( .A(cclow_cnt[8]), .B(n52), .Y(N33) );
endmodule


module SNPS_CLOCK_GATE_HIGH_updphy_FF_DEPTH_NUM34_FF_DEPTH_NBT6 ( CLK, EN, 
        ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module dbnc_WIDTH3 ( o_dbc, o_chg, i_org, clk, rstz );
  input i_org, clk, rstz;
  output o_dbc, o_chg;
  wire   d_org_0_, N14, N15, N16, N17, net10299, n4, n5, n6, n7, n8, n1, n2,
         n3;
  wire   [2:0] db_cnt;

  SNPS_CLOCK_GATE_HIGH_dbnc_WIDTH3 clk_gate_db_cnt_reg ( .CLK(clk), .EN(N14), 
        .ENCLK(net10299), .TE(1'b0) );
  DFFRQX1 d_org_reg_0_ ( .D(i_org), .C(clk), .XR(rstz), .Q(d_org_0_) );
  DFFRQX1 db_cnt_reg_2_ ( .D(N17), .C(net10299), .XR(rstz), .Q(db_cnt[2]) );
  DFFRQX1 db_cnt_reg_1_ ( .D(N16), .C(net10299), .XR(rstz), .Q(db_cnt[1]) );
  DFFRQX1 db_cnt_reg_0_ ( .D(N15), .C(net10299), .XR(rstz), .Q(db_cnt[0]) );
  DFFRQX1 d_org_reg_1_ ( .D(n8), .C(net10299), .XR(rstz), .Q(o_dbc) );
  NAND21X1 U3 ( .B(n5), .A(n4), .Y(n6) );
  OAI32X1 U4 ( .A(n6), .B(n1), .C(n2), .D(n6), .E(n3), .Y(N17) );
  NOR2X1 U5 ( .A(n7), .B(n6), .Y(N16) );
  XNOR2XL U6 ( .A(n2), .B(n1), .Y(n7) );
  NAND4X1 U7 ( .A(n5), .B(n1), .C(n2), .D(n3), .Y(N14) );
  XNOR2XL U8 ( .A(o_dbc), .B(d_org_0_), .Y(n5) );
  AO22AXL U9 ( .A(d_org_0_), .B(o_chg), .C(o_dbc), .D(o_chg), .Y(n8) );
  NOR2X1 U10 ( .A(n4), .B(n5), .Y(o_chg) );
  NAND3X1 U11 ( .A(db_cnt[1]), .B(db_cnt[0]), .C(db_cnt[2]), .Y(n4) );
  NOR2X1 U12 ( .A(db_cnt[0]), .B(n6), .Y(N15) );
  INVX1 U13 ( .A(db_cnt[0]), .Y(n1) );
  INVX1 U14 ( .A(db_cnt[1]), .Y(n2) );
  INVX1 U15 ( .A(db_cnt[2]), .Y(n3) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dbnc_WIDTH3 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module updprl_a0 ( r_spec, r_dat_spec, r_auto_txgdcrc, r_dat_portrole, 
        r_dat_datarole, r_auto_discard, r_set_cpmsgid, r_dat_cpmsgid, r_rdat, 
        r_rdy, pid_ccidle, r_discard, ptx_ack, ptx_txact, ptx_fifopop, 
        prx_fifopsh, prx_gdmsgrcvd, prx_eoprcvd, prx_rcvdords, prx_fifowdat, 
        pff_c0dat, prl_rdat, prl_txauto, prl_last, prl_txreq, prl_c0set, 
        prl_cany0, prl_cany0r, prl_cany0w, prl_idle, prl_discard, prl_GCTxDone, 
        prl_fsm, prl_cpmsgid, prl_cany0adr, clk, srstz );
  input [1:0] r_spec;
  input [1:0] r_dat_spec;
  input [2:0] r_dat_cpmsgid;
  input [7:0] r_rdat;
  input [2:0] prx_rcvdords;
  input [7:0] prx_fifowdat;
  input [47:0] pff_c0dat;
  output [7:0] prl_rdat;
  output [6:0] prl_txauto;
  output [3:0] prl_fsm;
  output [2:0] prl_cpmsgid;
  output [7:0] prl_cany0adr;
  input r_auto_txgdcrc, r_dat_portrole, r_dat_datarole, r_auto_discard,
         r_set_cpmsgid, r_rdy, pid_ccidle, r_discard, ptx_ack, ptx_txact,
         ptx_fifopop, prx_fifopsh, prx_gdmsgrcvd, prx_eoprcvd, clk, srstz;
  output prl_last, prl_txreq, prl_c0set, prl_cany0, prl_cany0r, prl_cany0w,
         prl_idle, prl_discard, prl_GCTxDone;
  wire   sendgdcrc, stoptimer, N40, N41, c0_iop, N113, N114, N115, N116, N117,
         N118, N119, N120, N135, N136, N137, N138, N139, N140, N141, N142,
         N143, N151, N152, N153, N154, N155, N156, N157, N158, N165, N166,
         N167, N168, N169, N170, N171, N172, N173, N189, N190, N191, N192,
         N193, N194, N196, N203, N204, N205, N206, net10322, net10328,
         net10333, net10338, net10343, n6, n8, n23, n26, n30, n36, n37, n38,
         n39, n62, n75, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n99, n100, n9, n10, n11, n12, n13, n17, n18,
         n19, n20, n21, n22, n24, n25, n27, n28, n29, n31, n32, n33, n34, n35,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n76, n93, n94, n95, n96, n97, n98, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129;
  wire   [1:0] PrlTo;
  wire   [8:0] c0_cnt;
  wire   [7:0] txbuf;

  PrlTimer_1112a0 u0_PrlTimer ( .to(PrlTo), .restart(sendgdcrc), .stop(
        stoptimer), .clk(clk), .srstz(n17) );
  SNPS_CLOCK_GATE_HIGH_updprl_a0_0 clk_gate_txbuf_reg ( .CLK(clk), .EN(N41), 
        .ENCLK(net10322), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_updprl_a0_4 clk_gate_c0_adr_reg ( .CLK(clk), .EN(N194), 
        .ENCLK(net10328), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_updprl_a0_3 clk_gate_cs_prcl_reg ( .CLK(clk), .EN(N189), 
        .ENCLK(net10333), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_updprl_a0_2 clk_gate_c0_cnt_reg ( .CLK(clk), .EN(N196), 
        .ENCLK(net10338), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_updprl_a0_1 clk_gate_CpMsgId_reg ( .CLK(clk), .EN(N203), 
        .ENCLK(net10343), .TE(1'b0) );
  updprl_a0_DW01_inc_0 r328 ( .A(prl_cany0adr), .SUM({N120, N119, N118, N117, 
        N116, N115, N114, N113}) );
  DFFQX1 c0_iop_reg ( .D(n99), .C(net10333), .Q(c0_iop) );
  DFFQX1 canyon_m0_reg ( .D(n100), .C(clk), .Q(prl_cany0) );
  DFFQX1 c0_adr_reg_2_ ( .D(N153), .C(net10328), .Q(prl_cany0adr[2]) );
  DFFQX1 c0_adr_reg_1_ ( .D(N152), .C(net10328), .Q(prl_cany0adr[1]) );
  DFFQX1 c0_adr_reg_3_ ( .D(N154), .C(net10328), .Q(prl_cany0adr[3]) );
  DFFQX1 c0_adr_reg_4_ ( .D(N155), .C(net10328), .Q(prl_cany0adr[4]) );
  DFFQX1 c0_adr_reg_5_ ( .D(N156), .C(net10328), .Q(prl_cany0adr[5]) );
  DFFQX1 c0_adr_reg_6_ ( .D(N157), .C(net10328), .Q(prl_cany0adr[6]) );
  DFFQX1 c0_adr_reg_0_ ( .D(N151), .C(net10328), .Q(prl_cany0adr[0]) );
  DFFQX1 c0_adr_reg_7_ ( .D(N158), .C(net10328), .Q(prl_cany0adr[7]) );
  DFFQX1 txbuf_reg_5_ ( .D(r_rdat[5]), .C(net10322), .Q(txbuf[5]) );
  DFFQX1 txbuf_reg_1_ ( .D(r_rdat[1]), .C(net10322), .Q(txbuf[1]) );
  DFFQX1 CpMsgId_reg_0_ ( .D(N204), .C(net10343), .Q(prl_cpmsgid[0]) );
  DFFQX1 txbuf_reg_3_ ( .D(r_rdat[3]), .C(net10322), .Q(txbuf[3]) );
  DFFQX1 txbuf_reg_4_ ( .D(r_rdat[4]), .C(net10322), .Q(txbuf[4]) );
  DFFQX1 CpMsgId_reg_2_ ( .D(N206), .C(net10343), .Q(prl_cpmsgid[2]) );
  DFFQX1 CpMsgId_reg_1_ ( .D(N205), .C(net10343), .Q(prl_cpmsgid[1]) );
  DFFQX1 c0_cnt_reg_4_ ( .D(N169), .C(net10338), .Q(c0_cnt[4]) );
  DFFQX1 c0_cnt_reg_5_ ( .D(N170), .C(net10338), .Q(c0_cnt[5]) );
  DFFQX1 c0_cnt_reg_1_ ( .D(N166), .C(net10338), .Q(c0_cnt[1]) );
  DFFQX1 c0_cnt_reg_3_ ( .D(N168), .C(net10338), .Q(c0_cnt[3]) );
  DFFQX1 txbuf_reg_0_ ( .D(r_rdat[0]), .C(net10322), .Q(txbuf[0]) );
  DFFQX1 c0_cnt_reg_2_ ( .D(N167), .C(net10338), .Q(c0_cnt[2]) );
  DFFQX1 c0_cnt_reg_8_ ( .D(N173), .C(net10338), .Q(c0_cnt[8]) );
  DFFQX1 c0_cnt_reg_7_ ( .D(N172), .C(net10338), .Q(c0_cnt[7]) );
  DFFQX1 c0_cnt_reg_6_ ( .D(N171), .C(net10338), .Q(c0_cnt[6]) );
  DFFQXL txbuf_reg_6_ ( .D(r_rdat[6]), .C(net10322), .Q(txbuf[6]) );
  DFFQXL txbuf_reg_2_ ( .D(r_rdat[2]), .C(net10322), .Q(txbuf[2]) );
  DFFQXL txbuf_reg_7_ ( .D(r_rdat[7]), .C(net10322), .Q(txbuf[7]) );
  DFFQX1 c0_cnt_reg_0_ ( .D(N165), .C(net10338), .Q(c0_cnt[0]) );
  DFFQX1 cs_prcl_reg_3_ ( .D(N193), .C(net10333), .Q(prl_fsm[3]) );
  DFFQX1 cs_prcl_reg_0_ ( .D(N190), .C(net10333), .Q(prl_fsm[0]) );
  DFFQX1 cs_prcl_reg_1_ ( .D(N191), .C(net10333), .Q(prl_fsm[1]) );
  DFFQX1 cs_prcl_reg_2_ ( .D(N192), .C(net10333), .Q(prl_fsm[2]) );
  INVX1 U3 ( .A(1'b0), .Y(prl_txauto[3]) );
  INVX1 U5 ( .A(1'b0), .Y(prl_txauto[5]) );
  INVX1 U7 ( .A(1'b1), .Y(prl_txauto[6]) );
  NAND21X1 U9 ( .B(n113), .A(n107), .Y(n105) );
  INVX1 U10 ( .A(n105), .Y(n112) );
  NAND21X1 U11 ( .B(prl_fsm[2]), .A(n29), .Y(n107) );
  INVX1 U12 ( .A(n28), .Y(n29) );
  INVX1 U13 ( .A(n110), .Y(n113) );
  INVX1 U14 ( .A(prl_fsm[3]), .Y(n27) );
  INVX1 U15 ( .A(n45), .Y(n9) );
  INVXL U16 ( .A(prl_fsm[0]), .Y(n43) );
  INVXL U17 ( .A(prl_fsm[1]), .Y(n32) );
  NAND32X1 U18 ( .B(prl_fsm[0]), .C(prl_fsm[2]), .A(n35), .Y(n98) );
  NAND21XL U19 ( .B(prl_fsm[0]), .A(prl_fsm[1]), .Y(n53) );
  AO22X1 U20 ( .A(txbuf[3]), .B(n112), .C(prl_cpmsgid[2]), .D(n108), .Y(
        prl_rdat[3]) );
  NAND32X1 U21 ( .B(n32), .C(n43), .A(n27), .Y(n28) );
  INVX1 U22 ( .A(n45), .Y(n59) );
  INVXL U23 ( .A(n33), .Y(n35) );
  NAND21X1 U24 ( .B(prl_fsm[3]), .A(n32), .Y(n33) );
  INVX2 U25 ( .A(n101), .Y(prl_cany0w) );
  INVX3 U26 ( .A(prx_fifopsh), .Y(n44) );
  NAND21X1 U27 ( .B(prl_txauto[4]), .A(ptx_fifopop), .Y(n46) );
  AO21XL U28 ( .B(n104), .C(n103), .A(n108), .Y(prl_last) );
  OAI22XL U29 ( .A(n112), .B(n31), .C(n126), .D(n96), .Y(n42) );
  AO21XL U30 ( .B(n98), .C(n110), .A(n18), .Y(n74) );
  NAND21XL U31 ( .B(n59), .A(n93), .Y(n55) );
  MUX2IXL U32 ( .D0(r_spec[0]), .D1(r_dat_spec[0]), .S(n12), .Y(n10) );
  AOI22XL U33 ( .A(n75), .B(n59), .C(n103), .D(ptx_ack), .Y(n22) );
  AO22AXL U34 ( .A(n49), .B(prx_fifopsh), .C(n50), .D(c0_iop), .Y(N194) );
  AO22XL U35 ( .A(n66), .B(prx_fifowdat[7]), .C(N142), .D(n59), .Y(N172) );
  AO22XL U36 ( .A(n66), .B(prx_fifowdat[6]), .C(N141), .D(n59), .Y(N171) );
  AO22XL U37 ( .A(n66), .B(n56), .C(N140), .D(n59), .Y(N170) );
  AO22XL U38 ( .A(n66), .B(prx_fifowdat[4]), .C(N139), .D(n59), .Y(N169) );
  AND2XL U39 ( .A(N143), .B(n9), .Y(N173) );
  OR2XL U40 ( .A(c0_cnt[7]), .B(n119), .Y(n120) );
  OR2XL U41 ( .A(n118), .B(c0_cnt[6]), .Y(n119) );
  OR2XL U42 ( .A(n117), .B(c0_cnt[5]), .Y(n118) );
  OR2XL U43 ( .A(n116), .B(c0_cnt[4]), .Y(n117) );
  OR2XL U44 ( .A(n115), .B(c0_cnt[3]), .Y(n116) );
  OR2XL U45 ( .A(n114), .B(c0_cnt[2]), .Y(n115) );
  OR2XL U46 ( .A(c0_cnt[1]), .B(c0_cnt[0]), .Y(n114) );
  AO22XL U47 ( .A(n66), .B(n57), .C(N138), .D(n59), .Y(N168) );
  AO22XL U48 ( .A(n66), .B(prx_fifowdat[2]), .C(N137), .D(n59), .Y(N167) );
  AO22XL U49 ( .A(n66), .B(n58), .C(N136), .D(n59), .Y(N166) );
  AO22XL U50 ( .A(n66), .B(n60), .C(N135), .D(n9), .Y(N165) );
  INVX1 U51 ( .A(r_discard), .Y(n69) );
  INVX1 U52 ( .A(n18), .Y(n17) );
  NOR21XL U53 ( .B(prx_gdmsgrcvd), .A(r_set_cpmsgid), .Y(n37) );
  NAND32X1 U54 ( .B(r_set_cpmsgid), .C(prx_gdmsgrcvd), .A(n17), .Y(N203) );
  INVX1 U55 ( .A(ptx_fifopop), .Y(n31) );
  INVX1 U56 ( .A(srstz), .Y(n18) );
  INVX1 U57 ( .A(n127), .Y(n57) );
  INVX1 U58 ( .A(prl_txauto[4]), .Y(n103) );
  INVX1 U59 ( .A(n23), .Y(prl_c0set) );
  INVX1 U60 ( .A(ptx_ack), .Y(n126) );
  INVX1 U61 ( .A(prx_fifowdat[3]), .Y(n127) );
  INVX1 U62 ( .A(n61), .Y(n64) );
  INVX1 U63 ( .A(n48), .Y(n54) );
  NAND21X1 U64 ( .B(n43), .A(n59), .Y(prl_txauto[4]) );
  NAND32X1 U65 ( .B(n45), .C(n44), .A(n43), .Y(n101) );
  INVXL U66 ( .A(n107), .Y(n108) );
  INVX1 U67 ( .A(n98), .Y(prl_idle) );
  OAI21X1 U68 ( .B(ptx_txact), .C(prl_txauto[4]), .A(n102), .Y(prl_txreq) );
  NAND31X1 U69 ( .C(prl_discard), .A(n8), .B(n69), .Y(n6) );
  NAND43X1 U70 ( .B(n94), .C(n42), .D(n41), .A(n40), .Y(N189) );
  OAI221X1 U71 ( .A(n122), .B(n67), .C(n98), .D(n34), .E(n47), .Y(n41) );
  OAI211X1 U72 ( .C(n73), .D(n18), .A(n72), .B(n71), .Y(N191) );
  AOI31XL U73 ( .A(n70), .B(n69), .C(n68), .D(n113), .Y(n73) );
  INVX1 U74 ( .A(n102), .Y(n68) );
  NAND4X1 U75 ( .A(n77), .B(n78), .C(n79), .D(n80), .Y(n23) );
  NOR4XL U76 ( .A(n84), .B(n85), .C(pff_c0dat[22]), .D(pff_c0dat[20]), .Y(n79)
         );
  NOR4XL U77 ( .A(n81), .B(n82), .C(pff_c0dat[36]), .D(pff_c0dat[34]), .Y(n80)
         );
  NOR42XL U78 ( .C(pff_c0dat[3]), .D(pff_c0dat[2]), .A(n90), .B(n91), .Y(n77)
         );
  NAND2X1 U79 ( .A(n39), .B(n17), .Y(N204) );
  AOI22X1 U80 ( .A(pff_c0dat[9]), .B(n37), .C(r_dat_cpmsgid[0]), .D(
        r_set_cpmsgid), .Y(n39) );
  NAND2X1 U81 ( .A(n38), .B(n17), .Y(N205) );
  AOI22X1 U82 ( .A(pff_c0dat[10]), .B(n37), .C(r_dat_cpmsgid[1]), .D(
        r_set_cpmsgid), .Y(n38) );
  NAND2X1 U83 ( .A(n36), .B(n17), .Y(N206) );
  AOI22X1 U84 ( .A(pff_c0dat[11]), .B(n37), .C(r_set_cpmsgid), .D(
        r_dat_cpmsgid[2]), .Y(n36) );
  INVX1 U85 ( .A(sendgdcrc), .Y(n34) );
  NAND42X1 U86 ( .C(n61), .D(n94), .A(n30), .B(n128), .Y(n72) );
  OAI211XL U87 ( .C(n18), .D(n107), .A(n76), .B(n71), .Y(N192) );
  OAI211X1 U88 ( .C(n94), .D(n93), .A(n76), .B(n74), .Y(N190) );
  INVX1 U89 ( .A(n63), .Y(n76) );
  OAI31XL U90 ( .A(n96), .B(n18), .C(n125), .D(n72), .Y(n63) );
  NAND21X1 U91 ( .B(n94), .A(n54), .Y(n71) );
  AOI21AX1 U92 ( .B(n125), .C(n23), .A(n95), .Y(n100) );
  INVX1 U93 ( .A(n94), .Y(n95) );
  AO22X1 U94 ( .A(N119), .B(n55), .C(n54), .D(prx_fifowdat[6]), .Y(N157) );
  AO22X1 U95 ( .A(N117), .B(n55), .C(n54), .D(prx_fifowdat[4]), .Y(N155) );
  INVX1 U96 ( .A(n124), .Y(n56) );
  INVXL U97 ( .A(prx_fifowdat[5]), .Y(n124) );
  AO22X1 U98 ( .A(N118), .B(n55), .C(n54), .D(n56), .Y(N156) );
  OR2X1 U99 ( .A(n8), .B(n67), .Y(n102) );
  AND3X1 U100 ( .A(n97), .B(n125), .C(ptx_ack), .Y(prl_GCTxDone) );
  INVX1 U101 ( .A(n96), .Y(n97) );
  INVX1 U102 ( .A(n70), .Y(prl_discard) );
  NAND21X1 U103 ( .B(n53), .A(n13), .Y(n61) );
  AO22X1 U104 ( .A(N116), .B(n55), .C(n54), .D(n57), .Y(N154) );
  NAND32X1 U105 ( .B(n43), .C(n52), .A(n35), .Y(n48) );
  AO22X1 U106 ( .A(N115), .B(n55), .C(n54), .D(prx_fifowdat[2]), .Y(N153) );
  AO22X1 U107 ( .A(N114), .B(n55), .C(n54), .D(n58), .Y(N152) );
  INVX1 U108 ( .A(n93), .Y(n66) );
  INVX1 U109 ( .A(n129), .Y(n58) );
  INVX1 U110 ( .A(n128), .Y(n60) );
  AO22AXL U111 ( .A(txbuf[6]), .B(n112), .C(n113), .D(n10), .Y(prl_rdat[6]) );
  AO21XL U112 ( .B(txbuf[5]), .C(n112), .A(n111), .Y(prl_rdat[5]) );
  NOR5X1 U113 ( .A(r_dat_datarole), .B(prx_rcvdords[2]), .C(prx_rcvdords[1]), 
        .D(n110), .E(n109), .Y(n111) );
  INVX1 U114 ( .A(prx_rcvdords[0]), .Y(n109) );
  AND2XL U115 ( .A(txbuf[4]), .B(n112), .Y(prl_rdat[4]) );
  AO22AXL U116 ( .A(txbuf[7]), .B(n112), .C(n113), .D(n11), .Y(prl_rdat[7]) );
  MUX2IX1 U117 ( .D0(r_spec[1]), .D1(r_dat_spec[1]), .S(n12), .Y(n11) );
  AO22XL U118 ( .A(txbuf[2]), .B(n112), .C(prl_cpmsgid[1]), .D(n108), .Y(
        prl_rdat[2]) );
  AO22XL U119 ( .A(txbuf[1]), .B(n112), .C(prl_cpmsgid[0]), .D(n108), .Y(
        prl_rdat[1]) );
  NAND32X1 U120 ( .B(prl_fsm[2]), .C(n53), .A(n27), .Y(n110) );
  NAND32XL U121 ( .B(prl_fsm[2]), .C(n27), .A(n32), .Y(n45) );
  OAI211XL U122 ( .C(r_dat_portrole), .D(n107), .A(n106), .B(n110), .Y(
        prl_rdat[0]) );
  NAND21XL U123 ( .B(n105), .A(txbuf[0]), .Y(n106) );
  AND2X1 U124 ( .A(r_spec[1]), .B(r_spec[0]), .Y(n12) );
  NOR4XL U125 ( .A(c0_cnt[6]), .B(c0_cnt[7]), .C(c0_cnt[8]), .D(n21), .Y(n104)
         );
  NAND42X1 U126 ( .C(c0_cnt[4]), .D(c0_cnt[5]), .A(n20), .B(n19), .Y(n21) );
  NOR2X1 U127 ( .A(c0_cnt[1]), .B(c0_cnt[0]), .Y(n20) );
  NOR2X1 U128 ( .A(c0_cnt[3]), .B(c0_cnt[2]), .Y(n19) );
  NAND21XL U129 ( .B(n28), .A(prl_fsm[2]), .Y(n93) );
  OAI21BX1 U130 ( .C(PrlTo[0]), .B(r_auto_discard), .A(n122), .Y(stoptimer) );
  INVX1 U131 ( .A(n6), .Y(n122) );
  NAND42X1 U132 ( .C(pff_c0dat[14]), .D(pff_c0dat[13]), .A(prx_gdmsgrcvd), .B(
        n89), .Y(n87) );
  NOR3XL U133 ( .A(pff_c0dat[15]), .B(pff_c0dat[18]), .C(pff_c0dat[16]), .Y(
        n89) );
  NAND21X1 U134 ( .B(r_rdy), .A(n51), .Y(N41) );
  NOR42XL U135 ( .C(pff_c0dat[24]), .D(pff_c0dat[21]), .A(n87), .B(n88), .Y(
        n78) );
  NAND3X1 U136 ( .A(pff_c0dat[17]), .B(pff_c0dat[12]), .C(pff_c0dat[19]), .Y(
        n88) );
  OAI21BBX1 U137 ( .A(r_auto_txgdcrc), .B(prx_gdmsgrcvd), .C(n23), .Y(
        sendgdcrc) );
  NAND32X1 U138 ( .B(n24), .C(n18), .A(n22), .Y(n94) );
  AND3XL U139 ( .A(N40), .B(prx_fifopsh), .C(n64), .Y(n24) );
  AOI21BBXL U140 ( .B(pid_ccidle), .C(prx_eoprcvd), .A(prl_fsm[0]), .Y(n75) );
  OA21X1 U141 ( .B(n66), .C(n65), .A(n95), .Y(N193) );
  AND3X1 U142 ( .A(prx_fifowdat[0]), .B(n30), .C(n64), .Y(n65) );
  ENOX1 U143 ( .A(n26), .B(n129), .C(n26), .D(c0_iop), .Y(n99) );
  NAND43X1 U144 ( .B(n53), .C(n94), .D(n52), .A(n30), .Y(n26) );
  INVX1 U145 ( .A(n71), .Y(n49) );
  NOR43XL U146 ( .B(n127), .C(n123), .D(n62), .A(prx_fifowdat[2]), .Y(n30) );
  NAND42X1 U147 ( .C(pff_c0dat[47]), .D(pff_c0dat[45]), .A(n125), .B(n83), .Y(
        n81) );
  NOR3XL U148 ( .A(pff_c0dat[42]), .B(pff_c0dat[44]), .C(pff_c0dat[43]), .Y(
        n83) );
  AND2X1 U149 ( .A(pff_c0dat[33]), .B(pff_c0dat[30]), .Y(n92) );
  NAND4X1 U150 ( .A(pff_c0dat[40]), .B(pff_c0dat[37]), .C(n92), .D(
        pff_c0dat[35]), .Y(n90) );
  NAND3X1 U151 ( .A(pff_c0dat[0]), .B(pff_c0dat[46]), .C(pff_c0dat[1]), .Y(n91) );
  AO22X1 U152 ( .A(N120), .B(n55), .C(n54), .D(prx_fifowdat[7]), .Y(N158) );
  OR3XL U153 ( .A(pff_c0dat[41]), .B(pff_c0dat[39]), .C(pff_c0dat[38]), .Y(n82) );
  OR3XL U154 ( .A(pff_c0dat[26]), .B(pff_c0dat[25]), .C(pff_c0dat[23]), .Y(n85) );
  NAND32X1 U155 ( .B(pff_c0dat[28]), .C(pff_c0dat[27]), .A(n86), .Y(n84) );
  NOR3XL U156 ( .A(pff_c0dat[29]), .B(pff_c0dat[32]), .C(pff_c0dat[31]), .Y(
        n86) );
  INVX1 U157 ( .A(prl_cany0), .Y(n125) );
  NAND2X1 U158 ( .A(pid_ccidle), .B(PrlTo[0]), .Y(n8) );
  NAND43X1 U159 ( .B(prl_fsm[1]), .C(prl_fsm[2]), .D(n43), .A(n27), .Y(n67) );
  NAND32X1 U160 ( .B(n25), .C(n67), .A(PrlTo[1]), .Y(n70) );
  INVX1 U161 ( .A(r_auto_discard), .Y(n25) );
  NAND32XL U162 ( .B(prl_fsm[1]), .C(prl_fsm[0]), .A(n13), .Y(n96) );
  AND2XL U163 ( .A(n27), .B(prl_fsm[2]), .Y(n13) );
  NAND21X1 U164 ( .B(n93), .A(pid_ccidle), .Y(n47) );
  AO22X1 U165 ( .A(N113), .B(n55), .C(n54), .D(n60), .Y(N151) );
  INVX1 U166 ( .A(prx_fifowdat[0]), .Y(n128) );
  INVXL U167 ( .A(prl_fsm[2]), .Y(n52) );
  INVX1 U168 ( .A(prx_fifowdat[1]), .Y(n129) );
  BUFX3 U169 ( .A(prx_rcvdords[2]), .Y(prl_txauto[2]) );
  BUFX3 U170 ( .A(prx_rcvdords[1]), .Y(prl_txauto[1]) );
  BUFX3 U171 ( .A(prx_rcvdords[0]), .Y(prl_txauto[0]) );
  AOI31XL U172 ( .A(n47), .B(n101), .C(n46), .D(n94), .Y(n50) );
  INVXL U173 ( .A(prl_cany0r), .Y(n51) );
  AND2XL U174 ( .A(n95), .B(prl_cany0r), .Y(N196) );
  OAI22X1 U175 ( .A(n44), .B(n93), .C(n104), .D(n46), .Y(prl_cany0r) );
  NOR3XL U176 ( .A(prx_fifowdat[5]), .B(prx_fifowdat[7]), .C(prx_fifowdat[6]), 
        .Y(n62) );
  INVXL U177 ( .A(prx_fifowdat[4]), .Y(n123) );
  AO21XL U178 ( .B(n48), .C(n61), .A(n44), .Y(n40) );
  INVX1 U179 ( .A(c0_cnt[0]), .Y(N135) );
  OAI21BBX1 U180 ( .A(c0_cnt[0]), .B(c0_cnt[1]), .C(n114), .Y(N136) );
  OAI21BBX1 U181 ( .A(n114), .B(c0_cnt[2]), .C(n115), .Y(N137) );
  OAI21BBX1 U182 ( .A(n115), .B(c0_cnt[3]), .C(n116), .Y(N138) );
  OAI21BBX1 U183 ( .A(n116), .B(c0_cnt[4]), .C(n117), .Y(N139) );
  OAI21BBX1 U184 ( .A(n117), .B(c0_cnt[5]), .C(n118), .Y(N140) );
  OAI21BBX1 U185 ( .A(n118), .B(c0_cnt[6]), .C(n119), .Y(N141) );
  XNOR2XL U186 ( .A(n119), .B(c0_cnt[7]), .Y(N142) );
  XNOR2XL U187 ( .A(c0_cnt[8]), .B(n120), .Y(N143) );
  NOR3XL U188 ( .A(prx_fifowdat[5]), .B(prx_fifowdat[7]), .C(prx_fifowdat[6]), 
        .Y(n121) );
  NAND43X1 U189 ( .B(prx_fifowdat[4]), .C(prx_fifowdat[3]), .D(prx_fifowdat[2]), .A(n121), .Y(N40) );
endmodule


module updprl_a0_DW01_inc_0 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  XOR2X1 U1 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_updprl_a0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_updprl_a0_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_updprl_a0_3 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_updprl_a0_4 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_updprl_a0_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module PrlTimer_1112a0 ( to, restart, stop, clk, srstz );
  output [1:0] to;
  input restart, stop, clk, srstz;
  wire   ena, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N18, N19,
         N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, net10360, n12,
         n1, n2, n3, n4, n5, n6, n7, n8, n9, n10;
  wire   [11:0] timer;

  SNPS_CLOCK_GATE_HIGH_PrlTimer_1112a0 clk_gate_timer_reg ( .CLK(clk), .EN(N18), .ENCLK(net10360), .TE(1'b0) );
  PrlTimer_1112a0_DW01_inc_0 add_25 ( .A(timer), .SUM({N15, N14, N13, N12, N11, 
        N10, N9, N8, N7, N6, N5, N4}) );
  DFFQX1 ena_reg ( .D(n12), .C(clk), .Q(ena) );
  DFFQX1 timer_reg_1_ ( .D(N20), .C(net10360), .Q(timer[1]) );
  DFFQX1 timer_reg_2_ ( .D(N21), .C(net10360), .Q(timer[2]) );
  DFFQX1 timer_reg_0_ ( .D(N19), .C(net10360), .Q(timer[0]) );
  DFFQX1 timer_reg_10_ ( .D(N29), .C(net10360), .Q(timer[10]) );
  DFFQX1 timer_reg_6_ ( .D(N25), .C(net10360), .Q(timer[6]) );
  DFFQX1 timer_reg_7_ ( .D(N26), .C(net10360), .Q(timer[7]) );
  DFFQX1 timer_reg_11_ ( .D(N30), .C(net10360), .Q(timer[11]) );
  DFFQX1 timer_reg_8_ ( .D(N27), .C(net10360), .Q(timer[8]) );
  DFFQX1 timer_reg_9_ ( .D(N28), .C(net10360), .Q(timer[9]) );
  DFFQX1 timer_reg_4_ ( .D(N23), .C(net10360), .Q(timer[4]) );
  DFFQX1 timer_reg_3_ ( .D(N22), .C(net10360), .Q(timer[3]) );
  DFFQX1 timer_reg_5_ ( .D(N24), .C(net10360), .Q(timer[5]) );
  BUFX3 U3 ( .A(n8), .Y(n1) );
  NAND3X1 U4 ( .A(srstz), .B(ena), .C(n9), .Y(n8) );
  INVX1 U5 ( .A(n2), .Y(to[0]) );
  AOI211X1 U6 ( .C(n3), .D(timer[9]), .A(timer[10]), .B(timer[11]), .Y(n2) );
  INVX1 U7 ( .A(n4), .Y(n3) );
  AOI211X1 U8 ( .C(timer[6]), .D(n5), .A(timer[8]), .B(timer[7]), .Y(n4) );
  AO21X1 U9 ( .B(timer[4]), .C(timer[3]), .A(timer[5]), .Y(n5) );
  INVX1 U10 ( .A(n6), .Y(n12) );
  AOI31X1 U11 ( .A(srstz), .B(n7), .C(ena), .D(restart), .Y(n6) );
  INVX1 U12 ( .A(stop), .Y(n7) );
  NOR21XL U13 ( .B(N15), .A(n1), .Y(N30) );
  NOR21XL U14 ( .B(N14), .A(n1), .Y(N29) );
  NOR21XL U15 ( .B(N13), .A(n1), .Y(N28) );
  NOR21XL U16 ( .B(N12), .A(n1), .Y(N27) );
  NOR21XL U17 ( .B(N11), .A(n8), .Y(N26) );
  NOR21XL U18 ( .B(N10), .A(n8), .Y(N25) );
  NOR21XL U19 ( .B(N9), .A(n8), .Y(N24) );
  NOR21XL U20 ( .B(N8), .A(n8), .Y(N23) );
  NOR21XL U21 ( .B(N7), .A(n8), .Y(N22) );
  NOR21XL U22 ( .B(N6), .A(n8), .Y(N21) );
  NOR21XL U23 ( .B(N5), .A(n8), .Y(N20) );
  NOR21XL U24 ( .B(N4), .A(n8), .Y(N19) );
  NAND31X1 U25 ( .C(restart), .A(n8), .B(srstz), .Y(N18) );
  NOR3XL U26 ( .A(to[1]), .B(stop), .C(restart), .Y(n9) );
  INVX1 U27 ( .A(n10), .Y(to[1]) );
  OAI31XL U28 ( .A(timer[10]), .B(timer[9]), .C(timer[8]), .D(timer[11]), .Y(
        n10) );
endmodule


module PrlTimer_1112a0_DW01_inc_0 ( A, SUM );
  input [11:0] A;
  output [11:0] SUM;

  wire   [11:2] carry;

  HAD1X1 U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .SO(SUM[10]) );
  HAD1X1 U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .SO(SUM[9]) );
  HAD1X1 U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .SO(SUM[8]) );
  HAD1X1 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .SO(SUM[7]) );
  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  XOR2X1 U1 ( .A(carry[11]), .B(A[11]), .Y(SUM[11]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_PrlTimer_1112a0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module phyff_DEPTH_NUM34_DEPTH_NBT6 ( r_psh, r_pop, prx_psh, ptx_pop, r_last, 
        r_unlock, i_lockena, r_fiforst, i_ccidle, r_wdat, prx_wdat, txreq, 
        ffack, rdat0, full, empty, one, half, obsd, dat_7_1, ptr, fifowdat, 
        fifopsh, clk, srstz );
  input [7:0] r_wdat;
  input [7:0] prx_wdat;
  output [1:0] ffack;
  output [7:0] rdat0;
  output [55:0] dat_7_1;
  output [5:0] ptr;
  output [7:0] fifowdat;
  input r_psh, r_pop, prx_psh, ptx_pop, r_last, r_unlock, i_lockena, r_fiforst,
         i_ccidle, clk, srstz;
  output txreq, full, empty, one, half, obsd, fifopsh;
  wire   ps_locked, locked, mem_8__7_, mem_8__6_, mem_8__5_, mem_8__4_,
         mem_8__3_, mem_8__2_, mem_8__1_, mem_8__0_, mem_9__7_, mem_9__6_,
         mem_9__5_, mem_9__4_, mem_9__3_, mem_9__2_, mem_9__1_, mem_9__0_,
         mem_10__7_, mem_10__6_, mem_10__5_, mem_10__4_, mem_10__3_,
         mem_10__2_, mem_10__1_, mem_10__0_, mem_11__7_, mem_11__6_,
         mem_11__5_, mem_11__4_, mem_11__3_, mem_11__2_, mem_11__1_,
         mem_11__0_, mem_12__7_, mem_12__6_, mem_12__5_, mem_12__4_,
         mem_12__3_, mem_12__2_, mem_12__1_, mem_12__0_, mem_13__7_,
         mem_13__6_, mem_13__5_, mem_13__4_, mem_13__3_, mem_13__2_,
         mem_13__1_, mem_13__0_, mem_14__7_, mem_14__6_, mem_14__5_,
         mem_14__4_, mem_14__3_, mem_14__2_, mem_14__1_, mem_14__0_,
         mem_15__7_, mem_15__6_, mem_15__5_, mem_15__4_, mem_15__3_,
         mem_15__2_, mem_15__1_, mem_15__0_, mem_16__7_, mem_16__6_,
         mem_16__5_, mem_16__4_, mem_16__3_, mem_16__2_, mem_16__1_,
         mem_16__0_, mem_17__7_, mem_17__6_, mem_17__5_, mem_17__4_,
         mem_17__3_, mem_17__2_, mem_17__1_, mem_17__0_, mem_18__7_,
         mem_18__6_, mem_18__5_, mem_18__4_, mem_18__3_, mem_18__2_,
         mem_18__1_, mem_18__0_, mem_19__7_, mem_19__6_, mem_19__5_,
         mem_19__4_, mem_19__3_, mem_19__2_, mem_19__1_, mem_19__0_,
         mem_20__7_, mem_20__6_, mem_20__5_, mem_20__4_, mem_20__3_,
         mem_20__2_, mem_20__1_, mem_20__0_, mem_21__7_, mem_21__6_,
         mem_21__5_, mem_21__4_, mem_21__3_, mem_21__2_, mem_21__1_,
         mem_21__0_, mem_22__7_, mem_22__6_, mem_22__5_, mem_22__4_,
         mem_22__3_, mem_22__2_, mem_22__1_, mem_22__0_, mem_23__7_,
         mem_23__6_, mem_23__5_, mem_23__4_, mem_23__3_, mem_23__2_,
         mem_23__1_, mem_23__0_, mem_24__7_, mem_24__6_, mem_24__5_,
         mem_24__4_, mem_24__3_, mem_24__2_, mem_24__1_, mem_24__0_,
         mem_25__7_, mem_25__6_, mem_25__5_, mem_25__4_, mem_25__3_,
         mem_25__2_, mem_25__1_, mem_25__0_, mem_26__7_, mem_26__6_,
         mem_26__5_, mem_26__4_, mem_26__3_, mem_26__2_, mem_26__1_,
         mem_26__0_, mem_27__7_, mem_27__6_, mem_27__5_, mem_27__4_,
         mem_27__3_, mem_27__2_, mem_27__1_, mem_27__0_, mem_28__7_,
         mem_28__6_, mem_28__5_, mem_28__4_, mem_28__3_, mem_28__2_,
         mem_28__1_, mem_28__0_, mem_29__7_, mem_29__6_, mem_29__5_,
         mem_29__4_, mem_29__3_, mem_29__2_, mem_29__1_, mem_29__0_,
         mem_30__7_, mem_30__6_, mem_30__5_, mem_30__4_, mem_30__3_,
         mem_30__2_, mem_30__1_, mem_30__0_, mem_31__7_, mem_31__6_,
         mem_31__5_, mem_31__4_, mem_31__3_, mem_31__2_, mem_31__1_,
         mem_31__0_, mem_32__7_, mem_32__6_, mem_32__5_, mem_32__4_,
         mem_32__3_, mem_32__2_, mem_32__1_, mem_32__0_, mem_33__7_,
         mem_33__6_, mem_33__5_, mem_33__4_, mem_33__3_, mem_33__2_,
         mem_33__1_, mem_33__0_, N693, N733, N734, N735, N736, N737, N738,
         N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749,
         N750, N751, N752, N753, N754, N755, N756, N757, N758, N759, N760,
         N761, N762, N763, N764, N765, N766, N767, N768, N769, N770, N771,
         N772, N773, N774, N775, N776, N777, N778, N779, N780, N781, N782,
         N783, N784, N785, N786, N787, N788, N789, N790, N791, N792, N793,
         N794, N795, N796, N797, N798, N799, N800, N801, N802, N803, N804,
         N805, N806, N807, N808, N809, N810, N811, N812, N813, N814, N815,
         N816, N817, N818, N819, N820, N821, N822, N823, N824, N825, N826,
         N827, N828, N829, N830, N831, N832, N833, N834, N835, N836, N837,
         N838, N839, N840, N841, N842, N843, N844, N845, N846, N847, N848,
         N849, N850, N851, N852, N853, N854, N855, N856, N857, N858, N859,
         N860, N861, N862, N863, N864, N865, N866, N867, N868, N869, N870,
         N871, N872, N873, N874, N875, N876, N877, N878, N879, N880, N881,
         N882, N883, N884, N885, N886, N887, N888, N889, N890, N891, N892,
         N893, N894, N895, N896, N897, N898, N899, N900, N901, N902, N903,
         N904, N905, N906, N907, N908, N909, N910, N911, N912, N913, N914,
         N915, N916, N917, N918, N919, N920, N921, N922, N923, N924, N925,
         N926, N927, N928, N929, N930, N931, N932, N933, N934, N935, N936,
         N937, N938, N939, N940, N941, N942, N943, N944, N945, N946, N947,
         N948, N949, N950, N951, N952, N953, N954, N955, N956, N957, N958,
         N959, N960, N961, N962, N963, N964, N965, N966, N967, N968, N969,
         N970, N971, N972, N973, N974, N975, N976, N977, N978, N979, N980,
         N981, N982, N983, N984, N985, N986, N987, N988, N989, N990, N991,
         N992, N993, N994, N995, N996, N997, N998, N999, N1000, N1001, N1002,
         N1003, N1004, N1005, N1006, N1007, N1008, N1009, N1010, N1011, N1012,
         N1013, N1014, N1015, N1016, N1017, N1018, N1019, N1020, N1021, N1022,
         N1023, N1024, N1025, N1026, N1027, N1028, N1029, N1030, N1035, N1036,
         N1037, N1038, N1039, N1040, N1041, N1042, N1043, N1044, N1045, N1046,
         N1053, N1054, N1055, N1056, N1057, N1058, N1059, N1157, N1159,
         net10378, net10384, net10389, net10394, net10399, net10404, net10409,
         net10414, net10419, net10424, net10429, net10434, net10439, net10444,
         net10449, net10454, net10459, net10464, net10469, net10474, net10479,
         net10484, net10489, net10494, net10499, net10504, net10509, net10514,
         net10519, net10524, net10529, net10534, net10539, net10544, net10549,
         gt_97_A_2_, gt_97_A_1_, gt_97_A_0_, add_101_B_0_, n1, n2, n3, n4, n5,
         n6, n7, n9, n10, n11, n13, n14, n15, n16, n17, n18, n19, n21, n22,
         n23, n24, n25, n26, n27, n29, n30, n31, n32, n33, n34, n35, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n54, n55, n56, n57, n58, n59, n60, n62, n63, n64, n65, n66, n67, n68,
         n70, n71, n72, n73, n74, n75, n76, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522;
  wire   [5:1] add_101_carry;
  wire   [5:1] sub_101_carry;

  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_0 clk_gate_mem_reg_0_ ( 
        .CLK(clk), .EN(N1022), .ENCLK(net10378), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_34 clk_gate_mem_reg_1_ ( 
        .CLK(clk), .EN(N1013), .ENCLK(net10384), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_33 clk_gate_mem_reg_2_ ( 
        .CLK(clk), .EN(N1004), .ENCLK(net10389), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_32 clk_gate_mem_reg_3_ ( 
        .CLK(clk), .EN(N995), .ENCLK(net10394), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_31 clk_gate_mem_reg_4_ ( 
        .CLK(clk), .EN(N986), .ENCLK(net10399), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_30 clk_gate_mem_reg_5_ ( 
        .CLK(clk), .EN(N977), .ENCLK(net10404), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_29 clk_gate_mem_reg_6_ ( 
        .CLK(clk), .EN(N968), .ENCLK(net10409), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_28 clk_gate_mem_reg_7_ ( 
        .CLK(clk), .EN(N959), .ENCLK(net10414), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_27 clk_gate_mem_reg_8_ ( 
        .CLK(clk), .EN(N950), .ENCLK(net10419), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_26 clk_gate_mem_reg_9_ ( 
        .CLK(clk), .EN(N941), .ENCLK(net10424), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_25 clk_gate_mem_reg_10_ ( 
        .CLK(clk), .EN(N932), .ENCLK(net10429), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_24 clk_gate_mem_reg_11_ ( 
        .CLK(clk), .EN(N923), .ENCLK(net10434), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_23 clk_gate_mem_reg_12_ ( 
        .CLK(clk), .EN(N914), .ENCLK(net10439), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_22 clk_gate_mem_reg_13_ ( 
        .CLK(clk), .EN(N905), .ENCLK(net10444), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_21 clk_gate_mem_reg_14_ ( 
        .CLK(clk), .EN(N896), .ENCLK(net10449), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_20 clk_gate_mem_reg_15_ ( 
        .CLK(clk), .EN(N887), .ENCLK(net10454), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_19 clk_gate_mem_reg_16_ ( 
        .CLK(clk), .EN(N878), .ENCLK(net10459), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_18 clk_gate_mem_reg_17_ ( 
        .CLK(clk), .EN(N869), .ENCLK(net10464), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_17 clk_gate_mem_reg_18_ ( 
        .CLK(clk), .EN(N860), .ENCLK(net10469), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_16 clk_gate_mem_reg_19_ ( 
        .CLK(clk), .EN(N851), .ENCLK(net10474), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_15 clk_gate_mem_reg_20_ ( 
        .CLK(clk), .EN(N842), .ENCLK(net10479), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_14 clk_gate_mem_reg_21_ ( 
        .CLK(clk), .EN(N833), .ENCLK(net10484), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_13 clk_gate_mem_reg_22_ ( 
        .CLK(clk), .EN(N824), .ENCLK(net10489), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_12 clk_gate_mem_reg_23_ ( 
        .CLK(clk), .EN(N815), .ENCLK(net10494), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_11 clk_gate_mem_reg_24_ ( 
        .CLK(clk), .EN(N806), .ENCLK(net10499), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_10 clk_gate_mem_reg_25_ ( 
        .CLK(clk), .EN(N797), .ENCLK(net10504), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_9 clk_gate_mem_reg_26_ ( 
        .CLK(clk), .EN(N788), .ENCLK(net10509), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_8 clk_gate_mem_reg_27_ ( 
        .CLK(clk), .EN(N779), .ENCLK(net10514), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_7 clk_gate_mem_reg_28_ ( 
        .CLK(clk), .EN(N770), .ENCLK(net10519), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_6 clk_gate_mem_reg_29_ ( 
        .CLK(clk), .EN(N761), .ENCLK(net10524), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_5 clk_gate_mem_reg_30_ ( 
        .CLK(clk), .EN(N752), .ENCLK(net10529), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_4 clk_gate_mem_reg_31_ ( 
        .CLK(clk), .EN(N743), .ENCLK(net10534), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_3 clk_gate_mem_reg_32_ ( 
        .CLK(clk), .EN(N734), .ENCLK(net10539), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_2 clk_gate_mem_reg_33_ ( 
        .CLK(clk), .EN(N733), .ENCLK(net10544), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_1 clk_gate_pshptr_reg ( 
        .CLK(clk), .EN(N1053), .ENCLK(net10549), .TE(1'b0) );
  DFFQX1 mem_reg_33__7_ ( .D(fifowdat[7]), .C(net10544), .Q(mem_33__7_) );
  DFFQX1 mem_reg_32__7_ ( .D(N742), .C(net10539), .Q(mem_32__7_) );
  DFFQX1 mem_reg_31__7_ ( .D(N751), .C(net10534), .Q(mem_31__7_) );
  DFFQX1 mem_reg_30__7_ ( .D(N760), .C(net10529), .Q(mem_30__7_) );
  DFFQX1 mem_reg_29__7_ ( .D(N769), .C(net10524), .Q(mem_29__7_) );
  DFFQX1 mem_reg_28__7_ ( .D(N778), .C(net10519), .Q(mem_28__7_) );
  DFFQX1 mem_reg_33__6_ ( .D(fifowdat[6]), .C(net10544), .Q(mem_33__6_) );
  DFFQX1 mem_reg_32__6_ ( .D(N741), .C(net10539), .Q(mem_32__6_) );
  DFFQX1 mem_reg_31__6_ ( .D(N750), .C(net10534), .Q(mem_31__6_) );
  DFFQX1 mem_reg_30__6_ ( .D(N759), .C(net10529), .Q(mem_30__6_) );
  DFFQX1 mem_reg_29__6_ ( .D(N768), .C(net10524), .Q(mem_29__6_) );
  DFFQX1 mem_reg_28__6_ ( .D(N777), .C(net10519), .Q(mem_28__6_) );
  DFFQX1 mem_reg_33__5_ ( .D(fifowdat[5]), .C(net10544), .Q(mem_33__5_) );
  DFFQX1 mem_reg_32__5_ ( .D(N740), .C(net10539), .Q(mem_32__5_) );
  DFFQX1 mem_reg_31__5_ ( .D(N749), .C(net10534), .Q(mem_31__5_) );
  DFFQX1 mem_reg_30__5_ ( .D(N758), .C(net10529), .Q(mem_30__5_) );
  DFFQX1 mem_reg_29__5_ ( .D(N767), .C(net10524), .Q(mem_29__5_) );
  DFFQX1 mem_reg_28__5_ ( .D(N776), .C(net10519), .Q(mem_28__5_) );
  DFFQX1 mem_reg_33__4_ ( .D(fifowdat[4]), .C(net10544), .Q(mem_33__4_) );
  DFFQX1 mem_reg_32__4_ ( .D(N739), .C(net10539), .Q(mem_32__4_) );
  DFFQX1 mem_reg_31__4_ ( .D(N748), .C(net10534), .Q(mem_31__4_) );
  DFFQX1 mem_reg_30__4_ ( .D(N757), .C(net10529), .Q(mem_30__4_) );
  DFFQX1 mem_reg_29__4_ ( .D(N766), .C(net10524), .Q(mem_29__4_) );
  DFFQX1 mem_reg_28__4_ ( .D(N775), .C(net10519), .Q(mem_28__4_) );
  DFFQX1 mem_reg_33__3_ ( .D(fifowdat[3]), .C(net10544), .Q(mem_33__3_) );
  DFFQX1 mem_reg_32__3_ ( .D(N738), .C(net10539), .Q(mem_32__3_) );
  DFFQX1 mem_reg_31__3_ ( .D(N747), .C(net10534), .Q(mem_31__3_) );
  DFFQX1 mem_reg_30__3_ ( .D(N756), .C(net10529), .Q(mem_30__3_) );
  DFFQX1 mem_reg_29__3_ ( .D(N765), .C(net10524), .Q(mem_29__3_) );
  DFFQX1 mem_reg_28__3_ ( .D(N774), .C(net10519), .Q(mem_28__3_) );
  DFFQX1 mem_reg_33__2_ ( .D(fifowdat[2]), .C(net10544), .Q(mem_33__2_) );
  DFFQX1 mem_reg_32__2_ ( .D(N737), .C(net10539), .Q(mem_32__2_) );
  DFFQX1 mem_reg_31__2_ ( .D(N746), .C(net10534), .Q(mem_31__2_) );
  DFFQX1 mem_reg_30__2_ ( .D(N755), .C(net10529), .Q(mem_30__2_) );
  DFFQX1 mem_reg_29__2_ ( .D(N764), .C(net10524), .Q(mem_29__2_) );
  DFFQX1 mem_reg_28__2_ ( .D(N773), .C(net10519), .Q(mem_28__2_) );
  DFFQX1 mem_reg_33__1_ ( .D(fifowdat[1]), .C(net10544), .Q(mem_33__1_) );
  DFFQX1 mem_reg_32__1_ ( .D(N736), .C(net10539), .Q(mem_32__1_) );
  DFFQX1 mem_reg_31__1_ ( .D(N745), .C(net10534), .Q(mem_31__1_) );
  DFFQX1 mem_reg_30__1_ ( .D(N754), .C(net10529), .Q(mem_30__1_) );
  DFFQX1 mem_reg_29__1_ ( .D(N763), .C(net10524), .Q(mem_29__1_) );
  DFFQX1 mem_reg_28__1_ ( .D(N772), .C(net10519), .Q(mem_28__1_) );
  DFFQX1 mem_reg_33__0_ ( .D(fifowdat[0]), .C(net10544), .Q(mem_33__0_) );
  DFFQX1 mem_reg_32__0_ ( .D(N735), .C(net10539), .Q(mem_32__0_) );
  DFFQX1 mem_reg_31__0_ ( .D(N744), .C(net10534), .Q(mem_31__0_) );
  DFFQX1 mem_reg_30__0_ ( .D(N753), .C(net10529), .Q(mem_30__0_) );
  DFFQX1 mem_reg_29__0_ ( .D(N762), .C(net10524), .Q(mem_29__0_) );
  DFFQX1 mem_reg_28__0_ ( .D(N771), .C(net10519), .Q(mem_28__0_) );
  DFFQX1 mem_reg_27__7_ ( .D(N787), .C(net10514), .Q(mem_27__7_) );
  DFFQX1 mem_reg_26__7_ ( .D(N796), .C(net10509), .Q(mem_26__7_) );
  DFFQX1 mem_reg_25__7_ ( .D(N805), .C(net10504), .Q(mem_25__7_) );
  DFFQX1 mem_reg_24__7_ ( .D(N814), .C(net10499), .Q(mem_24__7_) );
  DFFQX1 mem_reg_23__7_ ( .D(N823), .C(net10494), .Q(mem_23__7_) );
  DFFQX1 mem_reg_22__7_ ( .D(N832), .C(net10489), .Q(mem_22__7_) );
  DFFQX1 mem_reg_21__7_ ( .D(N841), .C(net10484), .Q(mem_21__7_) );
  DFFQX1 mem_reg_20__7_ ( .D(N850), .C(net10479), .Q(mem_20__7_) );
  DFFQX1 mem_reg_19__7_ ( .D(N859), .C(net10474), .Q(mem_19__7_) );
  DFFQX1 mem_reg_18__7_ ( .D(N868), .C(net10469), .Q(mem_18__7_) );
  DFFQX1 mem_reg_17__7_ ( .D(N877), .C(net10464), .Q(mem_17__7_) );
  DFFQX1 mem_reg_16__7_ ( .D(N886), .C(net10459), .Q(mem_16__7_) );
  DFFQX1 mem_reg_15__7_ ( .D(N895), .C(net10454), .Q(mem_15__7_) );
  DFFQX1 mem_reg_14__7_ ( .D(N904), .C(net10449), .Q(mem_14__7_) );
  DFFQX1 mem_reg_13__7_ ( .D(N913), .C(net10444), .Q(mem_13__7_) );
  DFFQX1 mem_reg_12__7_ ( .D(N922), .C(net10439), .Q(mem_12__7_) );
  DFFQX1 mem_reg_11__7_ ( .D(N931), .C(net10434), .Q(mem_11__7_) );
  DFFQX1 mem_reg_10__7_ ( .D(N940), .C(net10429), .Q(mem_10__7_) );
  DFFQX1 mem_reg_9__7_ ( .D(N949), .C(net10424), .Q(mem_9__7_) );
  DFFQX1 mem_reg_8__7_ ( .D(N958), .C(net10419), .Q(mem_8__7_) );
  DFFQX1 mem_reg_27__6_ ( .D(N786), .C(net10514), .Q(mem_27__6_) );
  DFFQX1 mem_reg_26__6_ ( .D(N795), .C(net10509), .Q(mem_26__6_) );
  DFFQX1 mem_reg_25__6_ ( .D(N804), .C(net10504), .Q(mem_25__6_) );
  DFFQX1 mem_reg_24__6_ ( .D(N813), .C(net10499), .Q(mem_24__6_) );
  DFFQX1 mem_reg_23__6_ ( .D(N822), .C(net10494), .Q(mem_23__6_) );
  DFFQX1 mem_reg_22__6_ ( .D(N831), .C(net10489), .Q(mem_22__6_) );
  DFFQX1 mem_reg_21__6_ ( .D(N840), .C(net10484), .Q(mem_21__6_) );
  DFFQX1 mem_reg_20__6_ ( .D(N849), .C(net10479), .Q(mem_20__6_) );
  DFFQX1 mem_reg_19__6_ ( .D(N858), .C(net10474), .Q(mem_19__6_) );
  DFFQX1 mem_reg_18__6_ ( .D(N867), .C(net10469), .Q(mem_18__6_) );
  DFFQX1 mem_reg_17__6_ ( .D(N876), .C(net10464), .Q(mem_17__6_) );
  DFFQX1 mem_reg_16__6_ ( .D(N885), .C(net10459), .Q(mem_16__6_) );
  DFFQX1 mem_reg_15__6_ ( .D(N894), .C(net10454), .Q(mem_15__6_) );
  DFFQX1 mem_reg_14__6_ ( .D(N903), .C(net10449), .Q(mem_14__6_) );
  DFFQX1 mem_reg_13__6_ ( .D(N912), .C(net10444), .Q(mem_13__6_) );
  DFFQX1 mem_reg_12__6_ ( .D(N921), .C(net10439), .Q(mem_12__6_) );
  DFFQX1 mem_reg_11__6_ ( .D(N930), .C(net10434), .Q(mem_11__6_) );
  DFFQX1 mem_reg_10__6_ ( .D(N939), .C(net10429), .Q(mem_10__6_) );
  DFFQX1 mem_reg_9__6_ ( .D(N948), .C(net10424), .Q(mem_9__6_) );
  DFFQX1 mem_reg_8__6_ ( .D(N957), .C(net10419), .Q(mem_8__6_) );
  DFFQX1 mem_reg_27__5_ ( .D(N785), .C(net10514), .Q(mem_27__5_) );
  DFFQX1 mem_reg_26__5_ ( .D(N794), .C(net10509), .Q(mem_26__5_) );
  DFFQX1 mem_reg_25__5_ ( .D(N803), .C(net10504), .Q(mem_25__5_) );
  DFFQX1 mem_reg_24__5_ ( .D(N812), .C(net10499), .Q(mem_24__5_) );
  DFFQX1 mem_reg_23__5_ ( .D(N821), .C(net10494), .Q(mem_23__5_) );
  DFFQX1 mem_reg_22__5_ ( .D(N830), .C(net10489), .Q(mem_22__5_) );
  DFFQX1 mem_reg_21__5_ ( .D(N839), .C(net10484), .Q(mem_21__5_) );
  DFFQX1 mem_reg_20__5_ ( .D(N848), .C(net10479), .Q(mem_20__5_) );
  DFFQX1 mem_reg_19__5_ ( .D(N857), .C(net10474), .Q(mem_19__5_) );
  DFFQX1 mem_reg_18__5_ ( .D(N866), .C(net10469), .Q(mem_18__5_) );
  DFFQX1 mem_reg_17__5_ ( .D(N875), .C(net10464), .Q(mem_17__5_) );
  DFFQX1 mem_reg_16__5_ ( .D(N884), .C(net10459), .Q(mem_16__5_) );
  DFFQX1 mem_reg_15__5_ ( .D(N893), .C(net10454), .Q(mem_15__5_) );
  DFFQX1 mem_reg_14__5_ ( .D(N902), .C(net10449), .Q(mem_14__5_) );
  DFFQX1 mem_reg_13__5_ ( .D(N911), .C(net10444), .Q(mem_13__5_) );
  DFFQX1 mem_reg_12__5_ ( .D(N920), .C(net10439), .Q(mem_12__5_) );
  DFFQX1 mem_reg_11__5_ ( .D(N929), .C(net10434), .Q(mem_11__5_) );
  DFFQX1 mem_reg_10__5_ ( .D(N938), .C(net10429), .Q(mem_10__5_) );
  DFFQX1 mem_reg_9__5_ ( .D(N947), .C(net10424), .Q(mem_9__5_) );
  DFFQX1 mem_reg_8__5_ ( .D(N956), .C(net10419), .Q(mem_8__5_) );
  DFFQX1 mem_reg_27__4_ ( .D(N784), .C(net10514), .Q(mem_27__4_) );
  DFFQX1 mem_reg_26__4_ ( .D(N793), .C(net10509), .Q(mem_26__4_) );
  DFFQX1 mem_reg_25__4_ ( .D(N802), .C(net10504), .Q(mem_25__4_) );
  DFFQX1 mem_reg_24__4_ ( .D(N811), .C(net10499), .Q(mem_24__4_) );
  DFFQX1 mem_reg_23__4_ ( .D(N820), .C(net10494), .Q(mem_23__4_) );
  DFFQX1 mem_reg_22__4_ ( .D(N829), .C(net10489), .Q(mem_22__4_) );
  DFFQX1 mem_reg_21__4_ ( .D(N838), .C(net10484), .Q(mem_21__4_) );
  DFFQX1 mem_reg_20__4_ ( .D(N847), .C(net10479), .Q(mem_20__4_) );
  DFFQX1 mem_reg_19__4_ ( .D(N856), .C(net10474), .Q(mem_19__4_) );
  DFFQX1 mem_reg_18__4_ ( .D(N865), .C(net10469), .Q(mem_18__4_) );
  DFFQX1 mem_reg_17__4_ ( .D(N874), .C(net10464), .Q(mem_17__4_) );
  DFFQX1 mem_reg_16__4_ ( .D(N883), .C(net10459), .Q(mem_16__4_) );
  DFFQX1 mem_reg_15__4_ ( .D(N892), .C(net10454), .Q(mem_15__4_) );
  DFFQX1 mem_reg_14__4_ ( .D(N901), .C(net10449), .Q(mem_14__4_) );
  DFFQX1 mem_reg_13__4_ ( .D(N910), .C(net10444), .Q(mem_13__4_) );
  DFFQX1 mem_reg_12__4_ ( .D(N919), .C(net10439), .Q(mem_12__4_) );
  DFFQX1 mem_reg_11__4_ ( .D(N928), .C(net10434), .Q(mem_11__4_) );
  DFFQX1 mem_reg_10__4_ ( .D(N937), .C(net10429), .Q(mem_10__4_) );
  DFFQX1 mem_reg_9__4_ ( .D(N946), .C(net10424), .Q(mem_9__4_) );
  DFFQX1 mem_reg_8__4_ ( .D(N955), .C(net10419), .Q(mem_8__4_) );
  DFFQX1 mem_reg_27__3_ ( .D(N783), .C(net10514), .Q(mem_27__3_) );
  DFFQX1 mem_reg_26__3_ ( .D(N792), .C(net10509), .Q(mem_26__3_) );
  DFFQX1 mem_reg_25__3_ ( .D(N801), .C(net10504), .Q(mem_25__3_) );
  DFFQX1 mem_reg_24__3_ ( .D(N810), .C(net10499), .Q(mem_24__3_) );
  DFFQX1 mem_reg_23__3_ ( .D(N819), .C(net10494), .Q(mem_23__3_) );
  DFFQX1 mem_reg_22__3_ ( .D(N828), .C(net10489), .Q(mem_22__3_) );
  DFFQX1 mem_reg_21__3_ ( .D(N837), .C(net10484), .Q(mem_21__3_) );
  DFFQX1 mem_reg_20__3_ ( .D(N846), .C(net10479), .Q(mem_20__3_) );
  DFFQX1 mem_reg_19__3_ ( .D(N855), .C(net10474), .Q(mem_19__3_) );
  DFFQX1 mem_reg_18__3_ ( .D(N864), .C(net10469), .Q(mem_18__3_) );
  DFFQX1 mem_reg_17__3_ ( .D(N873), .C(net10464), .Q(mem_17__3_) );
  DFFQX1 mem_reg_16__3_ ( .D(N882), .C(net10459), .Q(mem_16__3_) );
  DFFQX1 mem_reg_15__3_ ( .D(N891), .C(net10454), .Q(mem_15__3_) );
  DFFQX1 mem_reg_14__3_ ( .D(N900), .C(net10449), .Q(mem_14__3_) );
  DFFQX1 mem_reg_13__3_ ( .D(N909), .C(net10444), .Q(mem_13__3_) );
  DFFQX1 mem_reg_12__3_ ( .D(N918), .C(net10439), .Q(mem_12__3_) );
  DFFQX1 mem_reg_11__3_ ( .D(N927), .C(net10434), .Q(mem_11__3_) );
  DFFQX1 mem_reg_10__3_ ( .D(N936), .C(net10429), .Q(mem_10__3_) );
  DFFQX1 mem_reg_9__3_ ( .D(N945), .C(net10424), .Q(mem_9__3_) );
  DFFQX1 mem_reg_8__3_ ( .D(N954), .C(net10419), .Q(mem_8__3_) );
  DFFQX1 mem_reg_27__2_ ( .D(N782), .C(net10514), .Q(mem_27__2_) );
  DFFQX1 mem_reg_26__2_ ( .D(N791), .C(net10509), .Q(mem_26__2_) );
  DFFQX1 mem_reg_25__2_ ( .D(N800), .C(net10504), .Q(mem_25__2_) );
  DFFQX1 mem_reg_24__2_ ( .D(N809), .C(net10499), .Q(mem_24__2_) );
  DFFQX1 mem_reg_23__2_ ( .D(N818), .C(net10494), .Q(mem_23__2_) );
  DFFQX1 mem_reg_22__2_ ( .D(N827), .C(net10489), .Q(mem_22__2_) );
  DFFQX1 mem_reg_21__2_ ( .D(N836), .C(net10484), .Q(mem_21__2_) );
  DFFQX1 mem_reg_20__2_ ( .D(N845), .C(net10479), .Q(mem_20__2_) );
  DFFQX1 mem_reg_19__2_ ( .D(N854), .C(net10474), .Q(mem_19__2_) );
  DFFQX1 mem_reg_18__2_ ( .D(N863), .C(net10469), .Q(mem_18__2_) );
  DFFQX1 mem_reg_17__2_ ( .D(N872), .C(net10464), .Q(mem_17__2_) );
  DFFQX1 mem_reg_16__2_ ( .D(N881), .C(net10459), .Q(mem_16__2_) );
  DFFQX1 mem_reg_15__2_ ( .D(N890), .C(net10454), .Q(mem_15__2_) );
  DFFQX1 mem_reg_14__2_ ( .D(N899), .C(net10449), .Q(mem_14__2_) );
  DFFQX1 mem_reg_13__2_ ( .D(N908), .C(net10444), .Q(mem_13__2_) );
  DFFQX1 mem_reg_12__2_ ( .D(N917), .C(net10439), .Q(mem_12__2_) );
  DFFQX1 mem_reg_11__2_ ( .D(N926), .C(net10434), .Q(mem_11__2_) );
  DFFQX1 mem_reg_10__2_ ( .D(N935), .C(net10429), .Q(mem_10__2_) );
  DFFQX1 mem_reg_9__2_ ( .D(N944), .C(net10424), .Q(mem_9__2_) );
  DFFQX1 mem_reg_8__2_ ( .D(N953), .C(net10419), .Q(mem_8__2_) );
  DFFQX1 mem_reg_27__1_ ( .D(N781), .C(net10514), .Q(mem_27__1_) );
  DFFQX1 mem_reg_26__1_ ( .D(N790), .C(net10509), .Q(mem_26__1_) );
  DFFQX1 mem_reg_25__1_ ( .D(N799), .C(net10504), .Q(mem_25__1_) );
  DFFQX1 mem_reg_24__1_ ( .D(N808), .C(net10499), .Q(mem_24__1_) );
  DFFQX1 mem_reg_23__1_ ( .D(N817), .C(net10494), .Q(mem_23__1_) );
  DFFQX1 mem_reg_22__1_ ( .D(N826), .C(net10489), .Q(mem_22__1_) );
  DFFQX1 mem_reg_21__1_ ( .D(N835), .C(net10484), .Q(mem_21__1_) );
  DFFQX1 mem_reg_20__1_ ( .D(N844), .C(net10479), .Q(mem_20__1_) );
  DFFQX1 mem_reg_19__1_ ( .D(N853), .C(net10474), .Q(mem_19__1_) );
  DFFQX1 mem_reg_18__1_ ( .D(N862), .C(net10469), .Q(mem_18__1_) );
  DFFQX1 mem_reg_17__1_ ( .D(N871), .C(net10464), .Q(mem_17__1_) );
  DFFQX1 mem_reg_16__1_ ( .D(N880), .C(net10459), .Q(mem_16__1_) );
  DFFQX1 mem_reg_15__1_ ( .D(N889), .C(net10454), .Q(mem_15__1_) );
  DFFQX1 mem_reg_14__1_ ( .D(N898), .C(net10449), .Q(mem_14__1_) );
  DFFQX1 mem_reg_13__1_ ( .D(N907), .C(net10444), .Q(mem_13__1_) );
  DFFQX1 mem_reg_12__1_ ( .D(N916), .C(net10439), .Q(mem_12__1_) );
  DFFQX1 mem_reg_11__1_ ( .D(N925), .C(net10434), .Q(mem_11__1_) );
  DFFQX1 mem_reg_10__1_ ( .D(N934), .C(net10429), .Q(mem_10__1_) );
  DFFQX1 mem_reg_9__1_ ( .D(N943), .C(net10424), .Q(mem_9__1_) );
  DFFQX1 mem_reg_8__1_ ( .D(N952), .C(net10419), .Q(mem_8__1_) );
  DFFQX1 mem_reg_27__0_ ( .D(N780), .C(net10514), .Q(mem_27__0_) );
  DFFQX1 mem_reg_26__0_ ( .D(N789), .C(net10509), .Q(mem_26__0_) );
  DFFQX1 mem_reg_25__0_ ( .D(N798), .C(net10504), .Q(mem_25__0_) );
  DFFQX1 mem_reg_24__0_ ( .D(N807), .C(net10499), .Q(mem_24__0_) );
  DFFQX1 mem_reg_23__0_ ( .D(N816), .C(net10494), .Q(mem_23__0_) );
  DFFQX1 mem_reg_22__0_ ( .D(N825), .C(net10489), .Q(mem_22__0_) );
  DFFQX1 mem_reg_21__0_ ( .D(N834), .C(net10484), .Q(mem_21__0_) );
  DFFQX1 mem_reg_20__0_ ( .D(N843), .C(net10479), .Q(mem_20__0_) );
  DFFQX1 mem_reg_19__0_ ( .D(N852), .C(net10474), .Q(mem_19__0_) );
  DFFQX1 mem_reg_18__0_ ( .D(N861), .C(net10469), .Q(mem_18__0_) );
  DFFQX1 mem_reg_17__0_ ( .D(N870), .C(net10464), .Q(mem_17__0_) );
  DFFQX1 mem_reg_16__0_ ( .D(N879), .C(net10459), .Q(mem_16__0_) );
  DFFQX1 mem_reg_15__0_ ( .D(N888), .C(net10454), .Q(mem_15__0_) );
  DFFQX1 mem_reg_14__0_ ( .D(N897), .C(net10449), .Q(mem_14__0_) );
  DFFQX1 mem_reg_13__0_ ( .D(N906), .C(net10444), .Q(mem_13__0_) );
  DFFQX1 mem_reg_12__0_ ( .D(N915), .C(net10439), .Q(mem_12__0_) );
  DFFQX1 mem_reg_11__0_ ( .D(N924), .C(net10434), .Q(mem_11__0_) );
  DFFQX1 mem_reg_10__0_ ( .D(N933), .C(net10429), .Q(mem_10__0_) );
  DFFQX1 mem_reg_9__0_ ( .D(N942), .C(net10424), .Q(mem_9__0_) );
  DFFQX1 mem_reg_8__0_ ( .D(N951), .C(net10419), .Q(mem_8__0_) );
  DFFQX1 mem_reg_1__3_ ( .D(N1017), .C(net10384), .Q(dat_7_1[3]) );
  DFFQX1 mem_reg_1__2_ ( .D(N1016), .C(net10384), .Q(dat_7_1[2]) );
  DFFQX1 mem_reg_1__1_ ( .D(N1015), .C(net10384), .Q(dat_7_1[1]) );
  DFFQX1 mem_reg_1__0_ ( .D(N1014), .C(net10384), .Q(dat_7_1[0]) );
  DFFQX1 locked_reg ( .D(ps_locked), .C(clk), .Q(locked) );
  DFFQX1 mem_reg_7__7_ ( .D(N967), .C(net10414), .Q(dat_7_1[55]) );
  DFFQX1 mem_reg_6__7_ ( .D(N976), .C(net10409), .Q(dat_7_1[47]) );
  DFFQX1 mem_reg_7__6_ ( .D(N966), .C(net10414), .Q(dat_7_1[54]) );
  DFFQX1 mem_reg_6__6_ ( .D(N975), .C(net10409), .Q(dat_7_1[46]) );
  DFFQX1 mem_reg_7__5_ ( .D(N965), .C(net10414), .Q(dat_7_1[53]) );
  DFFQX1 mem_reg_6__5_ ( .D(N974), .C(net10409), .Q(dat_7_1[45]) );
  DFFQX1 mem_reg_6__4_ ( .D(N973), .C(net10409), .Q(dat_7_1[44]) );
  DFFQX1 mem_reg_7__3_ ( .D(N963), .C(net10414), .Q(dat_7_1[51]) );
  DFFQX1 mem_reg_6__3_ ( .D(N972), .C(net10409), .Q(dat_7_1[43]) );
  DFFQX1 mem_reg_6__2_ ( .D(N971), .C(net10409), .Q(dat_7_1[42]) );
  DFFQX1 mem_reg_7__1_ ( .D(N961), .C(net10414), .Q(dat_7_1[49]) );
  DFFQX1 mem_reg_7__0_ ( .D(N960), .C(net10414), .Q(dat_7_1[48]) );
  DFFQX1 mem_reg_6__0_ ( .D(N969), .C(net10409), .Q(dat_7_1[40]) );
  DFFQX1 mem_reg_5__7_ ( .D(N985), .C(net10404), .Q(dat_7_1[39]) );
  DFFQX1 mem_reg_4__7_ ( .D(N994), .C(net10399), .Q(dat_7_1[31]) );
  DFFQX1 mem_reg_4__6_ ( .D(N993), .C(net10399), .Q(dat_7_1[30]) );
  DFFQX1 mem_reg_5__5_ ( .D(N983), .C(net10404), .Q(dat_7_1[37]) );
  DFFQX1 mem_reg_4__5_ ( .D(N992), .C(net10399), .Q(dat_7_1[29]) );
  DFFQX1 mem_reg_4__4_ ( .D(N991), .C(net10399), .Q(dat_7_1[28]) );
  DFFQX1 mem_reg_4__3_ ( .D(N990), .C(net10399), .Q(dat_7_1[27]) );
  DFFQX1 mem_reg_4__2_ ( .D(N989), .C(net10399), .Q(dat_7_1[26]) );
  DFFQX1 mem_reg_5__1_ ( .D(N979), .C(net10404), .Q(dat_7_1[33]) );
  DFFQX1 mem_reg_5__0_ ( .D(N978), .C(net10404), .Q(dat_7_1[32]) );
  DFFQX1 mem_reg_4__0_ ( .D(N987), .C(net10399), .Q(dat_7_1[24]) );
  DFFQX1 mem_reg_3__3_ ( .D(N999), .C(net10394), .Q(dat_7_1[19]) );
  DFFQX1 mem_reg_3__2_ ( .D(N998), .C(net10394), .Q(dat_7_1[18]) );
  DFFQX1 mem_reg_3__1_ ( .D(N997), .C(net10394), .Q(dat_7_1[17]) );
  DFFQX1 mem_reg_3__0_ ( .D(N996), .C(net10394), .Q(dat_7_1[16]) );
  DFFQX1 mem_reg_2__7_ ( .D(N1012), .C(net10389), .Q(dat_7_1[15]) );
  DFFQX1 mem_reg_2__6_ ( .D(N1011), .C(net10389), .Q(dat_7_1[14]) );
  DFFQX1 mem_reg_2__5_ ( .D(N1010), .C(net10389), .Q(dat_7_1[13]) );
  DFFQX1 mem_reg_7__4_ ( .D(N964), .C(net10414), .Q(dat_7_1[52]) );
  DFFQX1 mem_reg_7__2_ ( .D(N962), .C(net10414), .Q(dat_7_1[50]) );
  DFFQX1 mem_reg_6__1_ ( .D(N970), .C(net10409), .Q(dat_7_1[41]) );
  DFFQX1 mem_reg_5__6_ ( .D(N984), .C(net10404), .Q(dat_7_1[38]) );
  DFFQX1 mem_reg_5__4_ ( .D(N982), .C(net10404), .Q(dat_7_1[36]) );
  DFFQX1 mem_reg_5__3_ ( .D(N981), .C(net10404), .Q(dat_7_1[35]) );
  DFFQX1 mem_reg_5__2_ ( .D(N980), .C(net10404), .Q(dat_7_1[34]) );
  DFFQX1 mem_reg_4__1_ ( .D(N988), .C(net10399), .Q(dat_7_1[25]) );
  DFFQX1 mem_reg_1__7_ ( .D(N1021), .C(net10384), .Q(dat_7_1[7]) );
  DFFQX1 mem_reg_1__6_ ( .D(N1020), .C(net10384), .Q(dat_7_1[6]) );
  DFFQX1 mem_reg_1__5_ ( .D(N1019), .C(net10384), .Q(dat_7_1[5]) );
  DFFQX1 mem_reg_1__4_ ( .D(N1018), .C(net10384), .Q(dat_7_1[4]) );
  DFFQX1 mem_reg_3__7_ ( .D(N1003), .C(net10394), .Q(dat_7_1[23]) );
  DFFQX1 mem_reg_3__6_ ( .D(N1002), .C(net10394), .Q(dat_7_1[22]) );
  DFFQX1 mem_reg_3__5_ ( .D(N1001), .C(net10394), .Q(dat_7_1[21]) );
  DFFQX1 mem_reg_3__4_ ( .D(N1000), .C(net10394), .Q(dat_7_1[20]) );
  DFFQX1 mem_reg_2__4_ ( .D(N1009), .C(net10389), .Q(dat_7_1[12]) );
  DFFQX1 mem_reg_2__3_ ( .D(N1008), .C(net10389), .Q(dat_7_1[11]) );
  DFFQX1 mem_reg_2__2_ ( .D(N1007), .C(net10389), .Q(dat_7_1[10]) );
  DFFQX1 mem_reg_2__1_ ( .D(N1006), .C(net10389), .Q(dat_7_1[9]) );
  DFFQX1 mem_reg_2__0_ ( .D(N1005), .C(net10389), .Q(dat_7_1[8]) );
  DFFQX1 mem_reg_0__5_ ( .D(N1028), .C(net10378), .Q(rdat0[5]) );
  DFFQX1 mem_reg_0__1_ ( .D(N1024), .C(net10378), .Q(rdat0[1]) );
  DFFQX1 mem_reg_0__7_ ( .D(N1030), .C(net10378), .Q(rdat0[7]) );
  DFFQX1 mem_reg_0__6_ ( .D(N1029), .C(net10378), .Q(rdat0[6]) );
  DFFQX1 mem_reg_0__4_ ( .D(N1027), .C(net10378), .Q(rdat0[4]) );
  DFFQX1 mem_reg_0__3_ ( .D(N1026), .C(net10378), .Q(rdat0[3]) );
  DFFQX1 mem_reg_0__2_ ( .D(N1025), .C(net10378), .Q(rdat0[2]) );
  DFFQX1 mem_reg_0__0_ ( .D(N1023), .C(net10378), .Q(rdat0[0]) );
  DFFQX1 pshptr_reg_5_ ( .D(N1059), .C(net10549), .Q(ptr[5]) );
  DFFQX1 pshptr_reg_1_ ( .D(N1055), .C(net10549), .Q(ptr[1]) );
  DFFQX1 pshptr_reg_3_ ( .D(N1057), .C(net10549), .Q(ptr[3]) );
  DFFQX1 pshptr_reg_2_ ( .D(N1056), .C(net10549), .Q(ptr[2]) );
  DFFQX1 pshptr_reg_0_ ( .D(N1054), .C(net10549), .Q(ptr[0]) );
  DFFQX1 pshptr_reg_4_ ( .D(N1058), .C(net10549), .Q(ptr[4]) );
  NAND2X1 U3 ( .A(n269), .B(n159), .Y(n1) );
  INVX1 U4 ( .A(n257), .Y(n2) );
  BUFX3 U5 ( .A(n376), .Y(n3) );
  BUFX3 U6 ( .A(n280), .Y(n4) );
  INVX1 U7 ( .A(gt_97_A_2_), .Y(n5) );
  BUFX3 U8 ( .A(n171), .Y(n6) );
  NOR3XL U9 ( .A(n87), .B(n86), .C(ptr[4]), .Y(one) );
  NAND32XL U10 ( .B(ptr[4]), .C(n87), .A(n86), .Y(n84) );
  NAND2XL U11 ( .A(ptr[5]), .B(n479), .Y(n365) );
  NAND2XL U12 ( .A(ptr[2]), .B(n479), .Y(n221) );
  NAND2XL U13 ( .A(ptr[1]), .B(n479), .Y(n283) );
  NAND2XL U14 ( .A(ptr[3]), .B(n479), .Y(n257) );
  NAND2XL U15 ( .A(ptr[4]), .B(n479), .Y(n318) );
  NAND2XL U16 ( .A(ptr[0]), .B(n479), .Y(n436) );
  INVX1 U17 ( .A(n16), .Y(n14) );
  INVX1 U18 ( .A(n16), .Y(n15) );
  INVX1 U19 ( .A(n16), .Y(n13) );
  INVX1 U20 ( .A(n96), .Y(n16) );
  INVX1 U21 ( .A(n81), .Y(n80) );
  INVX1 U22 ( .A(n81), .Y(n79) );
  INVX1 U23 ( .A(n73), .Y(n71) );
  INVX1 U24 ( .A(n73), .Y(n70) );
  INVX1 U25 ( .A(n65), .Y(n63) );
  INVX1 U26 ( .A(n65), .Y(n62) );
  INVX1 U27 ( .A(n57), .Y(n55) );
  INVX1 U28 ( .A(n57), .Y(n54) );
  INVX1 U29 ( .A(n73), .Y(n72) );
  INVX1 U30 ( .A(n65), .Y(n64) );
  INVX1 U31 ( .A(n57), .Y(n56) );
  INVX1 U32 ( .A(n49), .Y(n41) );
  INVX1 U33 ( .A(n40), .Y(n38) );
  INVX1 U34 ( .A(n32), .Y(n30) );
  INVX1 U35 ( .A(n24), .Y(n22) );
  INVX1 U36 ( .A(n40), .Y(n39) );
  INVX1 U37 ( .A(n32), .Y(n31) );
  INVX1 U38 ( .A(n24), .Y(n23) );
  INVX1 U39 ( .A(n81), .Y(n78) );
  INVX1 U40 ( .A(n125), .Y(n81) );
  INVX1 U41 ( .A(n48), .Y(n44) );
  INVX1 U42 ( .A(n48), .Y(n45) );
  INVX1 U43 ( .A(n48), .Y(n46) );
  INVX1 U44 ( .A(n48), .Y(n47) );
  INVX1 U45 ( .A(n122), .Y(n73) );
  INVX1 U46 ( .A(n119), .Y(n65) );
  INVX1 U47 ( .A(n115), .Y(n57) );
  INVX1 U48 ( .A(n48), .Y(n42) );
  INVX1 U49 ( .A(n48), .Y(n43) );
  INVX1 U50 ( .A(fifowdat[3]), .Y(n11) );
  INVX1 U51 ( .A(fifowdat[3]), .Y(n10) );
  INVX1 U52 ( .A(fifowdat[3]), .Y(n9) );
  NOR21XL U53 ( .B(n268), .A(n222), .Y(n258) );
  NOR21XL U54 ( .B(n364), .A(n319), .Y(n354) );
  AND2X1 U55 ( .A(n110), .B(n158), .Y(n148) );
  INVX1 U56 ( .A(n32), .Y(n29) );
  INVX1 U57 ( .A(n103), .Y(n32) );
  INVX1 U58 ( .A(n24), .Y(n21) );
  INVX1 U59 ( .A(n100), .Y(n24) );
  INVX1 U60 ( .A(n40), .Y(n37) );
  INVX1 U61 ( .A(n106), .Y(n40) );
  INVX1 U62 ( .A(n109), .Y(n49) );
  INVX1 U63 ( .A(n109), .Y(n48) );
  INVX1 U64 ( .A(fifowdat[4]), .Y(n76) );
  INVX1 U65 ( .A(fifowdat[4]), .Y(n75) );
  INVX1 U66 ( .A(fifowdat[5]), .Y(n68) );
  INVX1 U67 ( .A(fifowdat[5]), .Y(n67) );
  INVX1 U68 ( .A(fifowdat[6]), .Y(n60) );
  INVX1 U69 ( .A(fifowdat[6]), .Y(n59) );
  INVX1 U70 ( .A(fifowdat[7]), .Y(n52) );
  INVX1 U71 ( .A(fifowdat[7]), .Y(n51) );
  INVX1 U72 ( .A(fifowdat[4]), .Y(n74) );
  INVX1 U73 ( .A(fifowdat[5]), .Y(n66) );
  INVX1 U74 ( .A(fifowdat[6]), .Y(n58) );
  INVX1 U75 ( .A(fifowdat[7]), .Y(n50) );
  INVX1 U76 ( .A(n95), .Y(fifowdat[3]) );
  AOI21BBXL U77 ( .B(n183), .C(n280), .A(n281), .Y(n270) );
  AOI21BBXL U78 ( .B(n145), .C(n280), .A(n331), .Y(n332) );
  AOI21BBXL U79 ( .B(n130), .C(n280), .A(n330), .Y(n320) );
  AOI21BBXL U80 ( .B(n171), .C(n183), .A(n184), .Y(n173) );
  AOI21BBXL U81 ( .B(n111), .C(n280), .A(n306), .Y(n296) );
  AOI21BBXL U82 ( .B(n196), .C(n280), .A(n294), .Y(n284) );
  AOI21BBXL U83 ( .B(n132), .C(n280), .A(n317), .Y(n307) );
  AND2X1 U84 ( .A(n469), .B(n470), .Y(n459) );
  NAND3X1 U85 ( .A(n269), .B(n222), .C(N1159), .Y(n171) );
  NAND2X1 U86 ( .A(n269), .B(n159), .Y(n110) );
  AOI21BBXL U87 ( .B(n145), .C(n376), .A(n425), .Y(n426) );
  AOI21BBXL U88 ( .B(n145), .C(n171), .A(n234), .Y(n235) );
  AOI21BBXL U89 ( .B(n130), .C(n171), .A(n233), .Y(n223) );
  AOI21BBXL U90 ( .B(n130), .C(n376), .A(n424), .Y(n414) );
  AOI21BBXL U91 ( .B(n171), .C(n196), .A(n185), .Y(n186) );
  AOI21BBXL U92 ( .B(n171), .C(n172), .A(n159), .Y(n161) );
  AOI21BBXL U93 ( .B(n111), .C(n171), .A(n208), .Y(n198) );
  AOI21BBXL U94 ( .B(n111), .C(n376), .A(n401), .Y(n391) );
  AOI21BBXL U95 ( .B(n183), .C(n376), .A(n377), .Y(n366) );
  AOI21BBXL U96 ( .B(n196), .C(n376), .A(n389), .Y(n379) );
  AOI21BBXL U97 ( .B(n132), .C(n376), .A(n413), .Y(n403) );
  AOI21BBXL U98 ( .B(n110), .C(n132), .A(n108), .Y(n94) );
  AOI21BBXL U99 ( .B(n132), .C(n171), .A(n220), .Y(n210) );
  AOI21BBXL U100 ( .B(n1), .C(n145), .A(n133), .Y(n135) );
  AOI21BBXL U101 ( .B(n1), .C(n196), .A(n502), .Y(n492) );
  AOI21BBXL U102 ( .B(n110), .C(n183), .A(n490), .Y(n480) );
  AOI21BBXL U103 ( .B(n1), .C(n111), .A(n513), .Y(n503) );
  AOI21BBXL U104 ( .B(n110), .C(n130), .A(n131), .Y(n112) );
  AND2X1 U105 ( .A(n280), .B(n353), .Y(n343) );
  AND2X1 U106 ( .A(n171), .B(n256), .Y(n246) );
  AND2X1 U107 ( .A(n376), .B(n447), .Y(n437) );
  NAND21X1 U108 ( .B(empty), .A(n476), .Y(n109) );
  AO21X1 U109 ( .B(gt_97_A_0_), .C(empty), .A(n82), .Y(N1035) );
  INVX1 U110 ( .A(sub_101_carry[1]), .Y(n82) );
  INVX1 U111 ( .A(fifowdat[0]), .Y(n35) );
  INVX1 U112 ( .A(fifowdat[0]), .Y(n34) );
  INVX1 U113 ( .A(fifowdat[1]), .Y(n27) );
  INVX1 U114 ( .A(fifowdat[1]), .Y(n26) );
  INVX1 U115 ( .A(fifowdat[2]), .Y(n19) );
  INVX1 U116 ( .A(fifowdat[2]), .Y(n18) );
  INVX1 U117 ( .A(fifowdat[0]), .Y(n33) );
  INVX1 U118 ( .A(fifowdat[1]), .Y(n25) );
  INVX1 U119 ( .A(fifowdat[2]), .Y(n17) );
  INVX1 U120 ( .A(n123), .Y(fifowdat[4]) );
  INVX1 U121 ( .A(n117), .Y(fifowdat[6]) );
  INVX1 U122 ( .A(n120), .Y(fifowdat[5]) );
  INVX1 U123 ( .A(n113), .Y(fifowdat[7]) );
  AND3X1 U124 ( .A(ptr[4]), .B(ptr[0]), .C(n85), .Y(half) );
  NAND4X1 U125 ( .A(N1157), .B(n269), .C(n365), .D(n257), .Y(n280) );
  NOR21XL U126 ( .B(n458), .A(n365), .Y(n448) );
  NAND3X1 U127 ( .A(n269), .B(n365), .C(n378), .Y(n376) );
  INVX1 U128 ( .A(n257), .Y(N1159) );
  INVX1 U129 ( .A(n318), .Y(N1157) );
  NOR2X1 U130 ( .A(n7), .B(n90), .Y(ffack[0]) );
  AOI21X1 U131 ( .B(one), .C(r_pop), .A(n93), .Y(n7) );
  INVX1 U132 ( .A(n84), .Y(empty) );
  AO2222XL U133 ( .A(full), .B(r_psh), .C(r_pop), .D(empty), .E(n92), .F(n90), 
        .G(n89), .H(n93), .Y(ffack[1]) );
  NAND3X1 U134 ( .A(n283), .B(n221), .C(gt_97_A_0_), .Y(n183) );
  INVX1 U135 ( .A(n436), .Y(gt_97_A_0_) );
  NAND21X1 U136 ( .B(gt_97_A_0_), .A(n84), .Y(sub_101_carry[1]) );
  INVX1 U137 ( .A(n102), .Y(fifowdat[1]) );
  INVX1 U138 ( .A(n99), .Y(fifowdat[2]) );
  INVX1 U139 ( .A(n105), .Y(fifowdat[0]) );
  AND2X1 U140 ( .A(n84), .B(n83), .Y(obsd) );
  INVX1 U141 ( .A(srstz), .Y(n83) );
  INVX1 U142 ( .A(n87), .Y(n85) );
  OR4X1 U143 ( .A(ptr[5]), .B(ptr[1]), .C(ptr[2]), .D(ptr[3]), .Y(n87) );
  INVX1 U144 ( .A(ptr[0]), .Y(n86) );
  MUX2IXL U145 ( .D0(r_wdat[6]), .D1(prx_wdat[6]), .S(prx_psh), .Y(n117) );
  MUX2IXL U146 ( .D0(r_wdat[4]), .D1(prx_wdat[4]), .S(prx_psh), .Y(n123) );
  XOR2X1 U147 ( .A(N693), .B(add_101_carry[5]), .Y(N1046) );
  AND2X1 U148 ( .A(N1157), .B(add_101_carry[4]), .Y(add_101_carry[5]) );
  XOR2X1 U149 ( .A(add_101_carry[4]), .B(N1157), .Y(N1045) );
  AND2X1 U150 ( .A(N1159), .B(add_101_carry[3]), .Y(add_101_carry[4]) );
  XOR2X1 U151 ( .A(add_101_carry[3]), .B(n2), .Y(N1044) );
  AND2X1 U152 ( .A(gt_97_A_2_), .B(add_101_carry[2]), .Y(add_101_carry[3]) );
  XOR2X1 U153 ( .A(add_101_carry[2]), .B(gt_97_A_2_), .Y(N1043) );
  AND2X1 U154 ( .A(gt_97_A_1_), .B(add_101_carry[1]), .Y(add_101_carry[2]) );
  XOR2X1 U155 ( .A(add_101_carry[1]), .B(gt_97_A_1_), .Y(N1042) );
  XNOR2XL U156 ( .A(N693), .B(sub_101_carry[5]), .Y(N1040) );
  OR2X1 U157 ( .A(sub_101_carry[4]), .B(N1157), .Y(sub_101_carry[5]) );
  XNOR2XL U158 ( .A(sub_101_carry[4]), .B(N1157), .Y(N1039) );
  OR2X1 U159 ( .A(sub_101_carry[3]), .B(N1159), .Y(sub_101_carry[4]) );
  XNOR2XL U160 ( .A(sub_101_carry[3]), .B(n2), .Y(N1038) );
  OR2X1 U161 ( .A(sub_101_carry[2]), .B(gt_97_A_2_), .Y(sub_101_carry[3]) );
  XNOR2XL U162 ( .A(sub_101_carry[2]), .B(gt_97_A_2_), .Y(N1037) );
  OR2X1 U163 ( .A(sub_101_carry[1]), .B(gt_97_A_1_), .Y(sub_101_carry[2]) );
  XNOR2XL U164 ( .A(sub_101_carry[1]), .B(gt_97_A_1_), .Y(N1036) );
  AND2X1 U165 ( .A(add_101_B_0_), .B(gt_97_A_0_), .Y(add_101_carry[1]) );
  XOR2X1 U166 ( .A(gt_97_A_0_), .B(add_101_B_0_), .Y(N1041) );
  NOR4XL U167 ( .A(ptr[4]), .B(ptr[3]), .C(ptr[2]), .D(ptr[1]), .Y(n88) );
  NOR21XL U168 ( .B(ptr[5]), .A(n88), .Y(full) );
  NOR3XL U169 ( .A(n89), .B(n90), .C(n91), .Y(txreq) );
  INVX1 U170 ( .A(i_ccidle), .Y(n89) );
  INVX1 U171 ( .A(n91), .Y(n93) );
  NAND2X1 U172 ( .A(r_psh), .B(r_last), .Y(n91) );
  OAI211X1 U173 ( .C(n94), .D(n95), .A(n13), .B(n97), .Y(N999) );
  NAND2X1 U174 ( .A(dat_7_1[27]), .B(n98), .Y(n97) );
  OAI211X1 U175 ( .C(n94), .D(n99), .A(n21), .B(n101), .Y(N998) );
  NAND2X1 U176 ( .A(dat_7_1[26]), .B(n98), .Y(n101) );
  OAI211X1 U177 ( .C(n94), .D(n102), .A(n29), .B(n104), .Y(N997) );
  NAND2X1 U178 ( .A(dat_7_1[25]), .B(n98), .Y(n104) );
  OAI211X1 U179 ( .C(n94), .D(n105), .A(n37), .B(n107), .Y(N996) );
  NAND2X1 U180 ( .A(dat_7_1[24]), .B(n98), .Y(n107) );
  OAI22X1 U181 ( .A(n108), .B(n42), .C(n110), .D(n111), .Y(N995) );
  OAI211X1 U182 ( .C(n112), .D(n113), .A(n114), .B(n56), .Y(N994) );
  NAND2X1 U183 ( .A(dat_7_1[39]), .B(n116), .Y(n114) );
  OAI211X1 U184 ( .C(n112), .D(n117), .A(n118), .B(n64), .Y(N993) );
  NAND2X1 U185 ( .A(dat_7_1[38]), .B(n116), .Y(n118) );
  OAI211X1 U186 ( .C(n112), .D(n120), .A(n121), .B(n72), .Y(N992) );
  NAND2X1 U187 ( .A(dat_7_1[37]), .B(n116), .Y(n121) );
  OAI211X1 U188 ( .C(n112), .D(n123), .A(n124), .B(n125), .Y(N991) );
  NAND2X1 U189 ( .A(dat_7_1[36]), .B(n116), .Y(n124) );
  OAI211X1 U190 ( .C(n112), .D(n95), .A(n126), .B(n13), .Y(N990) );
  NAND2X1 U191 ( .A(dat_7_1[35]), .B(n116), .Y(n126) );
  OAI211X1 U192 ( .C(n112), .D(n99), .A(n127), .B(n21), .Y(N989) );
  NAND2X1 U193 ( .A(dat_7_1[34]), .B(n116), .Y(n127) );
  OAI211X1 U194 ( .C(n112), .D(n102), .A(n128), .B(n29), .Y(N988) );
  NAND2X1 U195 ( .A(dat_7_1[33]), .B(n116), .Y(n128) );
  OAI211X1 U196 ( .C(n112), .D(n105), .A(n129), .B(n37), .Y(N987) );
  NAND2X1 U197 ( .A(dat_7_1[32]), .B(n116), .Y(n129) );
  NOR21XL U198 ( .B(n112), .A(n44), .Y(n116) );
  OAI22X1 U199 ( .A(n1), .B(n132), .C(n131), .D(n42), .Y(N986) );
  NOR21XL U200 ( .B(n133), .A(n134), .Y(n131) );
  OAI211X1 U201 ( .C(n135), .D(n113), .A(n136), .B(n56), .Y(N985) );
  NAND2X1 U202 ( .A(dat_7_1[47]), .B(n137), .Y(n136) );
  OAI211X1 U203 ( .C(n135), .D(n117), .A(n138), .B(n64), .Y(N984) );
  NAND2X1 U204 ( .A(dat_7_1[46]), .B(n137), .Y(n138) );
  OAI211X1 U205 ( .C(n135), .D(n120), .A(n139), .B(n72), .Y(N983) );
  NAND2X1 U206 ( .A(dat_7_1[45]), .B(n137), .Y(n139) );
  OAI211X1 U207 ( .C(n135), .D(n123), .A(n140), .B(n125), .Y(N982) );
  NAND2X1 U208 ( .A(dat_7_1[44]), .B(n137), .Y(n140) );
  OAI211X1 U209 ( .C(n135), .D(n95), .A(n141), .B(n13), .Y(N981) );
  NAND2X1 U210 ( .A(dat_7_1[43]), .B(n137), .Y(n141) );
  OAI211X1 U211 ( .C(n135), .D(n99), .A(n142), .B(n21), .Y(N980) );
  NAND2X1 U212 ( .A(dat_7_1[42]), .B(n137), .Y(n142) );
  OAI211X1 U213 ( .C(n135), .D(n102), .A(n143), .B(n29), .Y(N979) );
  NAND2X1 U214 ( .A(dat_7_1[41]), .B(n137), .Y(n143) );
  OAI211X1 U215 ( .C(n135), .D(n105), .A(n144), .B(n37), .Y(N978) );
  NAND2X1 U216 ( .A(dat_7_1[40]), .B(n137), .Y(n144) );
  NOR21XL U217 ( .B(n135), .A(n44), .Y(n137) );
  OAI22X1 U218 ( .A(n110), .B(n130), .C(n133), .D(n42), .Y(N977) );
  NOR2X1 U219 ( .A(n146), .B(n147), .Y(n133) );
  OAI211X1 U220 ( .C(n148), .D(n113), .A(n149), .B(n56), .Y(N976) );
  NAND2X1 U221 ( .A(dat_7_1[55]), .B(n150), .Y(n149) );
  OAI211X1 U222 ( .C(n148), .D(n117), .A(n151), .B(n64), .Y(N975) );
  NAND2X1 U223 ( .A(dat_7_1[54]), .B(n150), .Y(n151) );
  OAI211X1 U224 ( .C(n148), .D(n120), .A(n152), .B(n72), .Y(N974) );
  NAND2X1 U225 ( .A(dat_7_1[53]), .B(n150), .Y(n152) );
  OAI211X1 U226 ( .C(n148), .D(n123), .A(n153), .B(n125), .Y(N973) );
  NAND2X1 U227 ( .A(dat_7_1[52]), .B(n150), .Y(n153) );
  OAI211X1 U228 ( .C(n148), .D(n11), .A(n154), .B(n13), .Y(N972) );
  NAND2X1 U229 ( .A(dat_7_1[51]), .B(n150), .Y(n154) );
  OAI211X1 U230 ( .C(n148), .D(n19), .A(n155), .B(n21), .Y(N971) );
  NAND2X1 U231 ( .A(dat_7_1[50]), .B(n150), .Y(n155) );
  OAI211X1 U232 ( .C(n148), .D(n27), .A(n156), .B(n29), .Y(N970) );
  NAND2X1 U233 ( .A(dat_7_1[49]), .B(n150), .Y(n156) );
  OAI211X1 U234 ( .C(n148), .D(n35), .A(n157), .B(n37), .Y(N969) );
  NAND2X1 U235 ( .A(dat_7_1[48]), .B(n150), .Y(n157) );
  NOR21XL U236 ( .B(n148), .A(n44), .Y(n150) );
  ENOX1 U237 ( .A(n110), .B(n145), .C(n158), .D(n48), .Y(N968) );
  NAND2X1 U238 ( .A(n159), .B(n160), .Y(n158) );
  OAI211X1 U239 ( .C(n161), .D(n52), .A(n162), .B(n55), .Y(N967) );
  NAND2X1 U240 ( .A(mem_8__7_), .B(n163), .Y(n162) );
  OAI211X1 U241 ( .C(n161), .D(n60), .A(n164), .B(n63), .Y(N966) );
  NAND2X1 U242 ( .A(mem_8__6_), .B(n163), .Y(n164) );
  OAI211X1 U243 ( .C(n161), .D(n68), .A(n165), .B(n71), .Y(N965) );
  NAND2X1 U244 ( .A(mem_8__5_), .B(n163), .Y(n165) );
  OAI211X1 U245 ( .C(n161), .D(n76), .A(n166), .B(n80), .Y(N964) );
  NAND2X1 U246 ( .A(mem_8__4_), .B(n163), .Y(n166) );
  OAI211X1 U247 ( .C(n161), .D(n11), .A(n167), .B(n13), .Y(N963) );
  NAND2X1 U248 ( .A(mem_8__3_), .B(n163), .Y(n167) );
  OAI211X1 U249 ( .C(n161), .D(n19), .A(n168), .B(n21), .Y(N962) );
  NAND2X1 U250 ( .A(mem_8__2_), .B(n163), .Y(n168) );
  OAI211X1 U251 ( .C(n161), .D(n27), .A(n169), .B(n29), .Y(N961) );
  NAND2X1 U252 ( .A(mem_8__1_), .B(n163), .Y(n169) );
  OAI211X1 U253 ( .C(n161), .D(n35), .A(n170), .B(n37), .Y(N960) );
  NAND2X1 U254 ( .A(mem_8__0_), .B(n163), .Y(n170) );
  NOR21XL U255 ( .B(n161), .A(n45), .Y(n163) );
  OAI22X1 U256 ( .A(n1), .B(n160), .C(n159), .D(n43), .Y(N959) );
  OAI211X1 U257 ( .C(n173), .D(n52), .A(n174), .B(n55), .Y(N958) );
  NAND2X1 U258 ( .A(mem_9__7_), .B(n175), .Y(n174) );
  OAI211X1 U259 ( .C(n173), .D(n60), .A(n176), .B(n63), .Y(N957) );
  NAND2X1 U260 ( .A(mem_9__6_), .B(n175), .Y(n176) );
  OAI211X1 U261 ( .C(n173), .D(n68), .A(n177), .B(n71), .Y(N956) );
  NAND2X1 U262 ( .A(mem_9__5_), .B(n175), .Y(n177) );
  OAI211X1 U263 ( .C(n173), .D(n76), .A(n178), .B(n80), .Y(N955) );
  NAND2X1 U264 ( .A(mem_9__4_), .B(n175), .Y(n178) );
  OAI211X1 U265 ( .C(n173), .D(n11), .A(n179), .B(n13), .Y(N954) );
  NAND2X1 U266 ( .A(mem_9__3_), .B(n175), .Y(n179) );
  OAI211X1 U267 ( .C(n173), .D(n19), .A(n180), .B(n21), .Y(N953) );
  NAND2X1 U268 ( .A(mem_9__2_), .B(n175), .Y(n180) );
  OAI211X1 U269 ( .C(n173), .D(n27), .A(n181), .B(n29), .Y(N952) );
  NAND2X1 U270 ( .A(mem_9__1_), .B(n175), .Y(n181) );
  OAI211X1 U271 ( .C(n173), .D(n35), .A(n182), .B(n37), .Y(N951) );
  NAND2X1 U272 ( .A(mem_9__0_), .B(n175), .Y(n182) );
  NOR21XL U273 ( .B(n173), .A(n45), .Y(n175) );
  OAI22X1 U274 ( .A(n6), .B(n172), .C(n184), .D(n43), .Y(N950) );
  AOI21AX1 U275 ( .B(gt_97_A_0_), .C(N1159), .A(n185), .Y(n184) );
  OAI211X1 U276 ( .C(n186), .D(n52), .A(n187), .B(n55), .Y(N949) );
  NAND2X1 U277 ( .A(mem_10__7_), .B(n188), .Y(n187) );
  OAI211X1 U278 ( .C(n186), .D(n60), .A(n189), .B(n63), .Y(N948) );
  NAND2X1 U279 ( .A(mem_10__6_), .B(n188), .Y(n189) );
  OAI211X1 U280 ( .C(n186), .D(n68), .A(n190), .B(n71), .Y(N947) );
  NAND2X1 U281 ( .A(mem_10__5_), .B(n188), .Y(n190) );
  OAI211X1 U282 ( .C(n186), .D(n76), .A(n191), .B(n80), .Y(N946) );
  NAND2X1 U283 ( .A(mem_10__4_), .B(n188), .Y(n191) );
  OAI211X1 U284 ( .C(n186), .D(n11), .A(n192), .B(n13), .Y(N945) );
  NAND2X1 U285 ( .A(mem_10__3_), .B(n188), .Y(n192) );
  OAI211X1 U286 ( .C(n186), .D(n19), .A(n193), .B(n21), .Y(N944) );
  NAND2X1 U287 ( .A(mem_10__2_), .B(n188), .Y(n193) );
  OAI211X1 U288 ( .C(n186), .D(n27), .A(n194), .B(n29), .Y(N943) );
  NAND2X1 U289 ( .A(mem_10__1_), .B(n188), .Y(n194) );
  OAI211X1 U290 ( .C(n186), .D(n35), .A(n195), .B(n37), .Y(N942) );
  NAND2X1 U291 ( .A(mem_10__0_), .B(n188), .Y(n195) );
  NOR21XL U292 ( .B(n186), .A(n45), .Y(n188) );
  OAI22X1 U293 ( .A(n6), .B(n183), .C(n185), .D(n43), .Y(N941) );
  AOI21X1 U294 ( .B(gt_97_A_1_), .C(N1159), .A(n197), .Y(n185) );
  OAI211X1 U295 ( .C(n198), .D(n52), .A(n199), .B(n55), .Y(N940) );
  NAND2X1 U296 ( .A(mem_11__7_), .B(n200), .Y(n199) );
  OAI211X1 U297 ( .C(n198), .D(n60), .A(n201), .B(n63), .Y(N939) );
  NAND2X1 U298 ( .A(mem_11__6_), .B(n200), .Y(n201) );
  OAI211X1 U299 ( .C(n198), .D(n68), .A(n202), .B(n71), .Y(N938) );
  NAND2X1 U300 ( .A(mem_11__5_), .B(n200), .Y(n202) );
  OAI211X1 U301 ( .C(n198), .D(n76), .A(n203), .B(n80), .Y(N937) );
  NAND2X1 U302 ( .A(mem_11__4_), .B(n200), .Y(n203) );
  OAI211X1 U303 ( .C(n198), .D(n11), .A(n204), .B(n13), .Y(N936) );
  NAND2X1 U304 ( .A(mem_11__3_), .B(n200), .Y(n204) );
  OAI211X1 U305 ( .C(n198), .D(n19), .A(n205), .B(n21), .Y(N935) );
  NAND2X1 U306 ( .A(mem_11__2_), .B(n200), .Y(n205) );
  OAI211X1 U307 ( .C(n198), .D(n27), .A(n206), .B(n29), .Y(N934) );
  NAND2X1 U308 ( .A(mem_11__1_), .B(n200), .Y(n206) );
  OAI211X1 U309 ( .C(n198), .D(n35), .A(n207), .B(n37), .Y(N933) );
  NAND2X1 U310 ( .A(mem_11__0_), .B(n200), .Y(n207) );
  NOR21XL U311 ( .B(n198), .A(n45), .Y(n200) );
  OAI22X1 U312 ( .A(n6), .B(n196), .C(n208), .D(n43), .Y(N932) );
  AOI21X1 U313 ( .B(n209), .C(N1159), .A(n197), .Y(n208) );
  OAI211X1 U314 ( .C(n210), .D(n52), .A(n211), .B(n55), .Y(N931) );
  NAND2X1 U315 ( .A(mem_12__7_), .B(n212), .Y(n211) );
  OAI211X1 U316 ( .C(n210), .D(n60), .A(n213), .B(n63), .Y(N930) );
  NAND2X1 U317 ( .A(mem_12__6_), .B(n212), .Y(n213) );
  OAI211X1 U318 ( .C(n210), .D(n68), .A(n214), .B(n71), .Y(N929) );
  NAND2X1 U319 ( .A(mem_12__5_), .B(n212), .Y(n214) );
  OAI211X1 U320 ( .C(n210), .D(n76), .A(n215), .B(n80), .Y(N928) );
  NAND2X1 U321 ( .A(mem_12__4_), .B(n212), .Y(n215) );
  OAI211X1 U322 ( .C(n210), .D(n11), .A(n216), .B(n14), .Y(N927) );
  NAND2X1 U323 ( .A(mem_12__3_), .B(n212), .Y(n216) );
  OAI211X1 U324 ( .C(n210), .D(n19), .A(n217), .B(n22), .Y(N926) );
  NAND2X1 U325 ( .A(mem_12__2_), .B(n212), .Y(n217) );
  OAI211X1 U326 ( .C(n210), .D(n27), .A(n218), .B(n30), .Y(N925) );
  NAND2X1 U327 ( .A(mem_12__1_), .B(n212), .Y(n218) );
  OAI211X1 U328 ( .C(n210), .D(n35), .A(n219), .B(n37), .Y(N924) );
  NAND2X1 U329 ( .A(mem_12__0_), .B(n212), .Y(n219) );
  NOR21XL U330 ( .B(n210), .A(n45), .Y(n212) );
  OAI22X1 U331 ( .A(n111), .B(n6), .C(n42), .D(n220), .Y(N923) );
  INVX1 U332 ( .A(n197), .Y(n220) );
  AOI21X1 U333 ( .B(n221), .C(n222), .A(n159), .Y(n197) );
  OAI211X1 U334 ( .C(n223), .D(n52), .A(n224), .B(n55), .Y(N922) );
  NAND2X1 U335 ( .A(mem_13__7_), .B(n225), .Y(n224) );
  OAI211X1 U336 ( .C(n223), .D(n60), .A(n226), .B(n63), .Y(N921) );
  NAND2X1 U337 ( .A(mem_13__6_), .B(n225), .Y(n226) );
  OAI211X1 U338 ( .C(n223), .D(n68), .A(n227), .B(n71), .Y(N920) );
  NAND2X1 U339 ( .A(mem_13__5_), .B(n225), .Y(n227) );
  OAI211X1 U340 ( .C(n223), .D(n76), .A(n228), .B(n80), .Y(N919) );
  NAND2X1 U341 ( .A(mem_13__4_), .B(n225), .Y(n228) );
  OAI211X1 U342 ( .C(n223), .D(n11), .A(n229), .B(n14), .Y(N918) );
  NAND2X1 U343 ( .A(mem_13__3_), .B(n225), .Y(n229) );
  OAI211X1 U344 ( .C(n223), .D(n19), .A(n230), .B(n22), .Y(N917) );
  NAND2X1 U345 ( .A(mem_13__2_), .B(n225), .Y(n230) );
  OAI211X1 U346 ( .C(n223), .D(n27), .A(n231), .B(n30), .Y(N916) );
  NAND2X1 U347 ( .A(mem_13__1_), .B(n225), .Y(n231) );
  OAI211X1 U348 ( .C(n223), .D(n35), .A(n232), .B(n37), .Y(N915) );
  NAND2X1 U349 ( .A(mem_13__0_), .B(n225), .Y(n232) );
  NOR21XL U350 ( .B(n223), .A(n45), .Y(n225) );
  OAI22X1 U351 ( .A(n132), .B(n6), .C(n233), .D(n43), .Y(N914) );
  AOI21AX1 U352 ( .B(n134), .C(N1159), .A(n234), .Y(n233) );
  OAI211X1 U353 ( .C(n235), .D(n52), .A(n236), .B(n55), .Y(N913) );
  NAND2X1 U354 ( .A(mem_14__7_), .B(n237), .Y(n236) );
  OAI211X1 U355 ( .C(n235), .D(n60), .A(n238), .B(n63), .Y(N912) );
  NAND2X1 U356 ( .A(mem_14__6_), .B(n237), .Y(n238) );
  OAI211X1 U357 ( .C(n235), .D(n68), .A(n239), .B(n71), .Y(N911) );
  NAND2X1 U358 ( .A(mem_14__5_), .B(n237), .Y(n239) );
  OAI211X1 U359 ( .C(n235), .D(n76), .A(n240), .B(n80), .Y(N910) );
  NAND2X1 U360 ( .A(mem_14__4_), .B(n237), .Y(n240) );
  OAI211X1 U361 ( .C(n235), .D(n11), .A(n241), .B(n14), .Y(N909) );
  NAND2X1 U362 ( .A(mem_14__3_), .B(n237), .Y(n241) );
  OAI211X1 U363 ( .C(n235), .D(n19), .A(n242), .B(n22), .Y(N908) );
  NAND2X1 U364 ( .A(mem_14__2_), .B(n237), .Y(n242) );
  OAI211X1 U365 ( .C(n235), .D(n27), .A(n243), .B(n30), .Y(N907) );
  NAND2X1 U366 ( .A(mem_14__1_), .B(n237), .Y(n243) );
  OAI211X1 U367 ( .C(n235), .D(n35), .A(n244), .B(n38), .Y(N906) );
  NAND2X1 U368 ( .A(mem_14__0_), .B(n237), .Y(n244) );
  NOR21XL U369 ( .B(n235), .A(n45), .Y(n237) );
  OAI22X1 U370 ( .A(n130), .B(n171), .C(n234), .D(n44), .Y(N905) );
  AOI21X1 U371 ( .B(n147), .C(N1159), .A(n245), .Y(n234) );
  OAI211X1 U372 ( .C(n246), .D(n52), .A(n247), .B(n55), .Y(N904) );
  NAND2X1 U373 ( .A(mem_15__7_), .B(n248), .Y(n247) );
  OAI211X1 U374 ( .C(n246), .D(n60), .A(n249), .B(n63), .Y(N903) );
  NAND2X1 U375 ( .A(mem_15__6_), .B(n248), .Y(n249) );
  OAI211X1 U376 ( .C(n246), .D(n68), .A(n250), .B(n71), .Y(N902) );
  NAND2X1 U377 ( .A(mem_15__5_), .B(n248), .Y(n250) );
  OAI211X1 U378 ( .C(n246), .D(n76), .A(n251), .B(n80), .Y(N901) );
  NAND2X1 U379 ( .A(mem_15__4_), .B(n248), .Y(n251) );
  OAI211X1 U380 ( .C(n246), .D(n11), .A(n252), .B(n14), .Y(N900) );
  NAND2X1 U381 ( .A(mem_15__3_), .B(n248), .Y(n252) );
  OAI211X1 U382 ( .C(n246), .D(n19), .A(n253), .B(n22), .Y(N899) );
  NAND2X1 U383 ( .A(mem_15__2_), .B(n248), .Y(n253) );
  OAI211X1 U384 ( .C(n246), .D(n27), .A(n254), .B(n30), .Y(N898) );
  NAND2X1 U385 ( .A(mem_15__1_), .B(n248), .Y(n254) );
  OAI211X1 U386 ( .C(n246), .D(n35), .A(n255), .B(n38), .Y(N897) );
  NAND2X1 U387 ( .A(mem_15__0_), .B(n248), .Y(n255) );
  NOR21XL U388 ( .B(n246), .A(n45), .Y(n248) );
  ENOX1 U389 ( .A(n145), .B(n6), .C(n256), .D(n48), .Y(N896) );
  OAI21X1 U390 ( .B(n257), .C(n160), .A(n222), .Y(n256) );
  OAI211X1 U391 ( .C(n258), .D(n52), .A(n259), .B(n55), .Y(N895) );
  NAND2X1 U392 ( .A(mem_16__7_), .B(n260), .Y(n259) );
  OAI211X1 U393 ( .C(n258), .D(n60), .A(n261), .B(n63), .Y(N894) );
  NAND2X1 U394 ( .A(mem_16__6_), .B(n260), .Y(n261) );
  OAI211X1 U395 ( .C(n258), .D(n68), .A(n262), .B(n71), .Y(N893) );
  NAND2X1 U396 ( .A(mem_16__5_), .B(n260), .Y(n262) );
  OAI211X1 U397 ( .C(n258), .D(n76), .A(n263), .B(n80), .Y(N892) );
  NAND2X1 U398 ( .A(mem_16__4_), .B(n260), .Y(n263) );
  OAI211X1 U399 ( .C(n258), .D(n11), .A(n264), .B(n14), .Y(N891) );
  NAND2X1 U400 ( .A(mem_16__3_), .B(n260), .Y(n264) );
  OAI211X1 U401 ( .C(n258), .D(n19), .A(n265), .B(n22), .Y(N890) );
  NAND2X1 U402 ( .A(mem_16__2_), .B(n260), .Y(n265) );
  OAI211X1 U403 ( .C(n258), .D(n27), .A(n266), .B(n30), .Y(N889) );
  NAND2X1 U404 ( .A(mem_16__1_), .B(n260), .Y(n266) );
  OAI211X1 U405 ( .C(n258), .D(n35), .A(n267), .B(n38), .Y(N888) );
  NAND2X1 U406 ( .A(mem_16__0_), .B(n260), .Y(n267) );
  NOR21XL U407 ( .B(n258), .A(n45), .Y(n260) );
  OAI22X1 U408 ( .A(n6), .B(n160), .C(n222), .D(n44), .Y(N887) );
  OAI211X1 U409 ( .C(n270), .D(n52), .A(n271), .B(n55), .Y(N886) );
  NAND2X1 U410 ( .A(mem_17__7_), .B(n272), .Y(n271) );
  OAI211X1 U411 ( .C(n270), .D(n60), .A(n273), .B(n63), .Y(N885) );
  NAND2X1 U412 ( .A(mem_17__6_), .B(n272), .Y(n273) );
  OAI211X1 U413 ( .C(n270), .D(n68), .A(n274), .B(n71), .Y(N884) );
  NAND2X1 U414 ( .A(mem_17__5_), .B(n272), .Y(n274) );
  OAI211X1 U415 ( .C(n270), .D(n76), .A(n275), .B(n80), .Y(N883) );
  NAND2X1 U416 ( .A(mem_17__4_), .B(n272), .Y(n275) );
  OAI211X1 U417 ( .C(n270), .D(n10), .A(n276), .B(n14), .Y(N882) );
  NAND2X1 U418 ( .A(mem_17__3_), .B(n272), .Y(n276) );
  OAI211X1 U419 ( .C(n270), .D(n18), .A(n277), .B(n22), .Y(N881) );
  NAND2X1 U420 ( .A(mem_17__2_), .B(n272), .Y(n277) );
  OAI211X1 U421 ( .C(n270), .D(n26), .A(n278), .B(n30), .Y(N880) );
  NAND2X1 U422 ( .A(mem_17__1_), .B(n272), .Y(n278) );
  OAI211X1 U423 ( .C(n270), .D(n34), .A(n279), .B(n38), .Y(N879) );
  NAND2X1 U424 ( .A(mem_17__0_), .B(n272), .Y(n279) );
  NOR21XL U425 ( .B(n270), .A(n45), .Y(n272) );
  OAI21X1 U426 ( .B(n41), .C(n281), .A(n268), .Y(N878) );
  OR2X1 U427 ( .A(n280), .B(n172), .Y(n268) );
  OAI31XL U428 ( .A(n282), .B(gt_97_A_0_), .C(N693), .D(n245), .Y(n281) );
  NAND3X1 U429 ( .A(n221), .B(n257), .C(n283), .Y(n282) );
  OAI211X1 U430 ( .C(n284), .D(n51), .A(n285), .B(n54), .Y(N877) );
  NAND2X1 U431 ( .A(mem_18__7_), .B(n286), .Y(n285) );
  OAI211X1 U432 ( .C(n284), .D(n59), .A(n287), .B(n62), .Y(N876) );
  NAND2X1 U433 ( .A(mem_18__6_), .B(n286), .Y(n287) );
  OAI211X1 U434 ( .C(n284), .D(n67), .A(n288), .B(n70), .Y(N875) );
  NAND2X1 U435 ( .A(mem_18__5_), .B(n286), .Y(n288) );
  OAI211X1 U436 ( .C(n284), .D(n75), .A(n289), .B(n79), .Y(N874) );
  NAND2X1 U437 ( .A(mem_18__4_), .B(n286), .Y(n289) );
  OAI211X1 U438 ( .C(n284), .D(n10), .A(n290), .B(n14), .Y(N873) );
  NAND2X1 U439 ( .A(mem_18__3_), .B(n286), .Y(n290) );
  OAI211X1 U440 ( .C(n284), .D(n18), .A(n291), .B(n22), .Y(N872) );
  NAND2X1 U441 ( .A(mem_18__2_), .B(n286), .Y(n291) );
  OAI211X1 U442 ( .C(n284), .D(n26), .A(n292), .B(n30), .Y(N871) );
  NAND2X1 U443 ( .A(mem_18__1_), .B(n286), .Y(n292) );
  OAI211X1 U444 ( .C(n284), .D(n34), .A(n293), .B(n38), .Y(N870) );
  NAND2X1 U445 ( .A(mem_18__0_), .B(n286), .Y(n293) );
  NOR21XL U446 ( .B(n284), .A(n46), .Y(n286) );
  OAI22X1 U447 ( .A(n183), .B(n4), .C(n294), .D(n44), .Y(N869) );
  AOI21X1 U448 ( .B(gt_97_A_1_), .C(N1157), .A(n295), .Y(n294) );
  OAI211X1 U449 ( .C(n296), .D(n51), .A(n297), .B(n54), .Y(N868) );
  NAND2X1 U450 ( .A(mem_19__7_), .B(n298), .Y(n297) );
  OAI211X1 U451 ( .C(n296), .D(n59), .A(n299), .B(n62), .Y(N867) );
  NAND2X1 U452 ( .A(mem_19__6_), .B(n298), .Y(n299) );
  OAI211X1 U453 ( .C(n296), .D(n67), .A(n300), .B(n70), .Y(N866) );
  NAND2X1 U454 ( .A(mem_19__5_), .B(n298), .Y(n300) );
  OAI211X1 U455 ( .C(n296), .D(n75), .A(n301), .B(n79), .Y(N865) );
  NAND2X1 U456 ( .A(mem_19__4_), .B(n298), .Y(n301) );
  OAI211X1 U457 ( .C(n296), .D(n10), .A(n302), .B(n14), .Y(N864) );
  NAND2X1 U458 ( .A(mem_19__3_), .B(n298), .Y(n302) );
  OAI211X1 U459 ( .C(n296), .D(n18), .A(n303), .B(n22), .Y(N863) );
  NAND2X1 U460 ( .A(mem_19__2_), .B(n298), .Y(n303) );
  OAI211X1 U461 ( .C(n296), .D(n26), .A(n304), .B(n30), .Y(N862) );
  NAND2X1 U462 ( .A(mem_19__1_), .B(n298), .Y(n304) );
  OAI211X1 U463 ( .C(n296), .D(n34), .A(n305), .B(n38), .Y(N861) );
  NAND2X1 U464 ( .A(mem_19__0_), .B(n298), .Y(n305) );
  NOR21XL U465 ( .B(n296), .A(n46), .Y(n298) );
  OAI22X1 U466 ( .A(n196), .B(n4), .C(n306), .D(n44), .Y(N860) );
  AOI21X1 U467 ( .B(n209), .C(N1157), .A(n295), .Y(n306) );
  OAI211X1 U468 ( .C(n307), .D(n51), .A(n308), .B(n54), .Y(N859) );
  NAND2X1 U469 ( .A(mem_20__7_), .B(n309), .Y(n308) );
  OAI211X1 U470 ( .C(n307), .D(n59), .A(n310), .B(n62), .Y(N858) );
  NAND2X1 U471 ( .A(mem_20__6_), .B(n309), .Y(n310) );
  OAI211X1 U472 ( .C(n307), .D(n67), .A(n311), .B(n70), .Y(N857) );
  NAND2X1 U473 ( .A(mem_20__5_), .B(n309), .Y(n311) );
  OAI211X1 U474 ( .C(n307), .D(n75), .A(n312), .B(n79), .Y(N856) );
  NAND2X1 U475 ( .A(mem_20__4_), .B(n309), .Y(n312) );
  OAI211X1 U476 ( .C(n307), .D(n10), .A(n313), .B(n14), .Y(N855) );
  NAND2X1 U477 ( .A(mem_20__3_), .B(n309), .Y(n313) );
  OAI211X1 U478 ( .C(n307), .D(n18), .A(n314), .B(n22), .Y(N854) );
  NAND2X1 U479 ( .A(mem_20__2_), .B(n309), .Y(n314) );
  OAI211X1 U480 ( .C(n307), .D(n26), .A(n315), .B(n30), .Y(N853) );
  NAND2X1 U481 ( .A(mem_20__1_), .B(n309), .Y(n315) );
  OAI211X1 U482 ( .C(n307), .D(n34), .A(n316), .B(n38), .Y(N852) );
  NAND2X1 U483 ( .A(mem_20__0_), .B(n309), .Y(n316) );
  NOR21XL U484 ( .B(n307), .A(n46), .Y(n309) );
  OAI22X1 U485 ( .A(n111), .B(n4), .C(n317), .D(n44), .Y(N851) );
  INVX1 U486 ( .A(n295), .Y(n317) );
  OAI21X1 U487 ( .B(n221), .C(n318), .A(n319), .Y(n295) );
  OAI211X1 U488 ( .C(n320), .D(n51), .A(n321), .B(n54), .Y(N850) );
  NAND2X1 U489 ( .A(mem_21__7_), .B(n322), .Y(n321) );
  OAI211X1 U490 ( .C(n320), .D(n59), .A(n323), .B(n62), .Y(N849) );
  NAND2X1 U491 ( .A(mem_21__6_), .B(n322), .Y(n323) );
  OAI211X1 U492 ( .C(n320), .D(n67), .A(n324), .B(n70), .Y(N848) );
  NAND2X1 U493 ( .A(mem_21__5_), .B(n322), .Y(n324) );
  OAI211X1 U494 ( .C(n320), .D(n75), .A(n325), .B(n79), .Y(N847) );
  NAND2X1 U495 ( .A(mem_21__4_), .B(n322), .Y(n325) );
  OAI211X1 U496 ( .C(n320), .D(n10), .A(n326), .B(n14), .Y(N846) );
  NAND2X1 U497 ( .A(mem_21__3_), .B(n322), .Y(n326) );
  OAI211X1 U498 ( .C(n320), .D(n18), .A(n327), .B(n22), .Y(N845) );
  NAND2X1 U499 ( .A(mem_21__2_), .B(n322), .Y(n327) );
  OAI211X1 U500 ( .C(n320), .D(n26), .A(n328), .B(n30), .Y(N844) );
  NAND2X1 U501 ( .A(mem_21__1_), .B(n322), .Y(n328) );
  OAI211X1 U502 ( .C(n320), .D(n34), .A(n329), .B(n38), .Y(N843) );
  NAND2X1 U503 ( .A(mem_21__0_), .B(n322), .Y(n329) );
  NOR21XL U504 ( .B(n320), .A(n46), .Y(n322) );
  OAI22X1 U505 ( .A(n132), .B(n4), .C(n330), .D(n44), .Y(N842) );
  AOI21AX1 U506 ( .B(n134), .C(N1157), .A(n331), .Y(n330) );
  OAI211X1 U507 ( .C(n332), .D(n51), .A(n333), .B(n54), .Y(N841) );
  NAND2X1 U508 ( .A(mem_22__7_), .B(n334), .Y(n333) );
  OAI211X1 U509 ( .C(n332), .D(n59), .A(n335), .B(n62), .Y(N840) );
  NAND2X1 U510 ( .A(mem_22__6_), .B(n334), .Y(n335) );
  OAI211X1 U511 ( .C(n332), .D(n67), .A(n336), .B(n70), .Y(N839) );
  NAND2X1 U512 ( .A(mem_22__5_), .B(n334), .Y(n336) );
  OAI211X1 U513 ( .C(n332), .D(n75), .A(n337), .B(n79), .Y(N838) );
  NAND2X1 U514 ( .A(mem_22__4_), .B(n334), .Y(n337) );
  OAI211X1 U515 ( .C(n332), .D(n10), .A(n338), .B(n15), .Y(N837) );
  NAND2X1 U516 ( .A(mem_22__3_), .B(n334), .Y(n338) );
  OAI211X1 U517 ( .C(n332), .D(n18), .A(n339), .B(n23), .Y(N836) );
  NAND2X1 U518 ( .A(mem_22__2_), .B(n334), .Y(n339) );
  OAI211X1 U519 ( .C(n332), .D(n26), .A(n340), .B(n31), .Y(N835) );
  NAND2X1 U520 ( .A(mem_22__1_), .B(n334), .Y(n340) );
  OAI211X1 U521 ( .C(n332), .D(n34), .A(n341), .B(n38), .Y(N834) );
  NAND2X1 U522 ( .A(mem_22__0_), .B(n334), .Y(n341) );
  NOR21XL U523 ( .B(n332), .A(n46), .Y(n334) );
  OAI22X1 U524 ( .A(n130), .B(n4), .C(n331), .D(n43), .Y(N833) );
  AOI21X1 U525 ( .B(n147), .C(N1157), .A(n342), .Y(n331) );
  OAI211X1 U526 ( .C(n343), .D(n51), .A(n344), .B(n54), .Y(N832) );
  NAND2X1 U527 ( .A(mem_23__7_), .B(n345), .Y(n344) );
  OAI211X1 U528 ( .C(n343), .D(n59), .A(n346), .B(n62), .Y(N831) );
  NAND2X1 U529 ( .A(mem_23__6_), .B(n345), .Y(n346) );
  OAI211X1 U530 ( .C(n343), .D(n67), .A(n347), .B(n70), .Y(N830) );
  NAND2X1 U531 ( .A(mem_23__5_), .B(n345), .Y(n347) );
  OAI211X1 U532 ( .C(n343), .D(n75), .A(n348), .B(n79), .Y(N829) );
  NAND2X1 U533 ( .A(mem_23__4_), .B(n345), .Y(n348) );
  OAI211X1 U534 ( .C(n343), .D(n10), .A(n349), .B(n15), .Y(N828) );
  NAND2X1 U535 ( .A(mem_23__3_), .B(n345), .Y(n349) );
  OAI211X1 U536 ( .C(n343), .D(n18), .A(n350), .B(n23), .Y(N827) );
  NAND2X1 U537 ( .A(mem_23__2_), .B(n345), .Y(n350) );
  OAI211X1 U538 ( .C(n343), .D(n26), .A(n351), .B(n31), .Y(N826) );
  NAND2X1 U539 ( .A(mem_23__1_), .B(n345), .Y(n351) );
  OAI211X1 U540 ( .C(n343), .D(n34), .A(n352), .B(n38), .Y(N825) );
  NAND2X1 U541 ( .A(mem_23__0_), .B(n345), .Y(n352) );
  NOR21XL U542 ( .B(n343), .A(n46), .Y(n345) );
  ENOX1 U543 ( .A(n145), .B(n4), .C(n353), .D(n49), .Y(N824) );
  OAI21X1 U544 ( .B(n160), .C(n318), .A(n319), .Y(n353) );
  OAI211X1 U545 ( .C(n354), .D(n51), .A(n355), .B(n54), .Y(N823) );
  NAND2X1 U546 ( .A(mem_24__7_), .B(n356), .Y(n355) );
  OAI211X1 U547 ( .C(n354), .D(n59), .A(n357), .B(n62), .Y(N822) );
  NAND2X1 U548 ( .A(mem_24__6_), .B(n356), .Y(n357) );
  OAI211X1 U549 ( .C(n354), .D(n67), .A(n358), .B(n70), .Y(N821) );
  NAND2X1 U550 ( .A(mem_24__5_), .B(n356), .Y(n358) );
  OAI211X1 U551 ( .C(n354), .D(n75), .A(n359), .B(n79), .Y(N820) );
  NAND2X1 U552 ( .A(mem_24__4_), .B(n356), .Y(n359) );
  OAI211X1 U553 ( .C(n354), .D(n10), .A(n360), .B(n15), .Y(N819) );
  NAND2X1 U554 ( .A(mem_24__3_), .B(n356), .Y(n360) );
  OAI211X1 U555 ( .C(n354), .D(n18), .A(n361), .B(n23), .Y(N818) );
  NAND2X1 U556 ( .A(mem_24__2_), .B(n356), .Y(n361) );
  OAI211X1 U557 ( .C(n354), .D(n26), .A(n362), .B(n31), .Y(N817) );
  NAND2X1 U558 ( .A(mem_24__1_), .B(n356), .Y(n362) );
  OAI211X1 U559 ( .C(n354), .D(n34), .A(n363), .B(n39), .Y(N816) );
  NAND2X1 U560 ( .A(mem_24__0_), .B(n356), .Y(n363) );
  NOR21XL U561 ( .B(n354), .A(n46), .Y(n356) );
  OAI22X1 U562 ( .A(n160), .B(n280), .C(n319), .D(n43), .Y(N815) );
  INVX1 U563 ( .A(n342), .Y(n319) );
  OAI211X1 U564 ( .C(n366), .D(n51), .A(n367), .B(n54), .Y(N814) );
  NAND2X1 U565 ( .A(mem_25__7_), .B(n368), .Y(n367) );
  OAI211X1 U566 ( .C(n366), .D(n59), .A(n369), .B(n62), .Y(N813) );
  NAND2X1 U567 ( .A(mem_25__6_), .B(n368), .Y(n369) );
  OAI211X1 U568 ( .C(n366), .D(n67), .A(n370), .B(n70), .Y(N812) );
  NAND2X1 U569 ( .A(mem_25__5_), .B(n368), .Y(n370) );
  OAI211X1 U570 ( .C(n366), .D(n75), .A(n371), .B(n79), .Y(N811) );
  NAND2X1 U571 ( .A(mem_25__4_), .B(n368), .Y(n371) );
  OAI211X1 U572 ( .C(n366), .D(n10), .A(n372), .B(n15), .Y(N810) );
  NAND2X1 U573 ( .A(mem_25__3_), .B(n368), .Y(n372) );
  OAI211X1 U574 ( .C(n366), .D(n18), .A(n373), .B(n23), .Y(N809) );
  NAND2X1 U575 ( .A(mem_25__2_), .B(n368), .Y(n373) );
  OAI211X1 U576 ( .C(n366), .D(n26), .A(n374), .B(n31), .Y(N808) );
  NAND2X1 U577 ( .A(mem_25__1_), .B(n368), .Y(n374) );
  OAI211X1 U578 ( .C(n366), .D(n34), .A(n375), .B(n39), .Y(N807) );
  NAND2X1 U579 ( .A(mem_25__0_), .B(n368), .Y(n375) );
  NOR21XL U580 ( .B(n366), .A(n46), .Y(n368) );
  OAI21X1 U581 ( .B(n377), .C(n41), .A(n364), .Y(N806) );
  OR2X1 U582 ( .A(n376), .B(n172), .Y(n364) );
  AOI21X1 U583 ( .B(n172), .C(n378), .A(N693), .Y(n377) );
  OAI211X1 U584 ( .C(n379), .D(n51), .A(n380), .B(n54), .Y(N805) );
  NAND2X1 U585 ( .A(mem_26__7_), .B(n381), .Y(n380) );
  OAI211X1 U586 ( .C(n379), .D(n59), .A(n382), .B(n62), .Y(N804) );
  NAND2X1 U587 ( .A(mem_26__6_), .B(n381), .Y(n382) );
  OAI211X1 U588 ( .C(n379), .D(n67), .A(n383), .B(n70), .Y(N803) );
  NAND2X1 U589 ( .A(mem_26__5_), .B(n381), .Y(n383) );
  OAI211X1 U590 ( .C(n379), .D(n75), .A(n384), .B(n79), .Y(N802) );
  NAND2X1 U591 ( .A(mem_26__4_), .B(n381), .Y(n384) );
  OAI211X1 U592 ( .C(n379), .D(n10), .A(n385), .B(n15), .Y(N801) );
  NAND2X1 U593 ( .A(mem_26__3_), .B(n381), .Y(n385) );
  OAI211X1 U594 ( .C(n379), .D(n18), .A(n386), .B(n23), .Y(N800) );
  NAND2X1 U595 ( .A(mem_26__2_), .B(n381), .Y(n386) );
  OAI211X1 U596 ( .C(n379), .D(n26), .A(n387), .B(n31), .Y(N799) );
  NAND2X1 U597 ( .A(mem_26__1_), .B(n381), .Y(n387) );
  OAI211X1 U598 ( .C(n379), .D(n34), .A(n388), .B(n39), .Y(N798) );
  NAND2X1 U599 ( .A(mem_26__0_), .B(n381), .Y(n388) );
  NOR21XL U600 ( .B(n379), .A(n46), .Y(n381) );
  OAI22X1 U601 ( .A(n183), .B(n3), .C(n389), .D(n43), .Y(N797) );
  AOI21X1 U602 ( .B(gt_97_A_1_), .C(n378), .A(n390), .Y(n389) );
  OAI211X1 U603 ( .C(n391), .D(n51), .A(n392), .B(n54), .Y(N796) );
  NAND2X1 U604 ( .A(mem_27__7_), .B(n393), .Y(n392) );
  OAI211X1 U605 ( .C(n391), .D(n59), .A(n394), .B(n62), .Y(N795) );
  NAND2X1 U606 ( .A(mem_27__6_), .B(n393), .Y(n394) );
  OAI211X1 U607 ( .C(n391), .D(n67), .A(n395), .B(n70), .Y(N794) );
  NAND2X1 U608 ( .A(mem_27__5_), .B(n393), .Y(n395) );
  OAI211X1 U609 ( .C(n391), .D(n75), .A(n396), .B(n79), .Y(N793) );
  NAND2X1 U610 ( .A(mem_27__4_), .B(n393), .Y(n396) );
  OAI211X1 U611 ( .C(n391), .D(n9), .A(n397), .B(n15), .Y(N792) );
  NAND2X1 U612 ( .A(mem_27__3_), .B(n393), .Y(n397) );
  OAI211X1 U613 ( .C(n391), .D(n17), .A(n398), .B(n23), .Y(N791) );
  NAND2X1 U614 ( .A(mem_27__2_), .B(n393), .Y(n398) );
  OAI211X1 U615 ( .C(n391), .D(n25), .A(n399), .B(n31), .Y(N790) );
  NAND2X1 U616 ( .A(mem_27__1_), .B(n393), .Y(n399) );
  OAI211X1 U617 ( .C(n391), .D(n33), .A(n400), .B(n39), .Y(N789) );
  NAND2X1 U618 ( .A(mem_27__0_), .B(n393), .Y(n400) );
  NOR21XL U619 ( .B(n391), .A(n46), .Y(n393) );
  OAI22X1 U620 ( .A(n196), .B(n3), .C(n401), .D(n43), .Y(N788) );
  AOI21X1 U621 ( .B(n209), .C(n378), .A(n390), .Y(n401) );
  OAI21X1 U622 ( .B(n221), .C(n402), .A(n365), .Y(n390) );
  OAI211X1 U623 ( .C(n403), .D(n50), .A(n404), .B(n56), .Y(N787) );
  NAND2X1 U624 ( .A(mem_28__7_), .B(n405), .Y(n404) );
  OAI211X1 U625 ( .C(n403), .D(n58), .A(n406), .B(n64), .Y(N786) );
  NAND2X1 U626 ( .A(mem_28__6_), .B(n405), .Y(n406) );
  OAI211X1 U627 ( .C(n403), .D(n66), .A(n407), .B(n72), .Y(N785) );
  NAND2X1 U628 ( .A(mem_28__5_), .B(n405), .Y(n407) );
  OAI211X1 U629 ( .C(n403), .D(n74), .A(n408), .B(n78), .Y(N784) );
  NAND2X1 U630 ( .A(mem_28__4_), .B(n405), .Y(n408) );
  OAI211X1 U631 ( .C(n403), .D(n9), .A(n409), .B(n15), .Y(N783) );
  NAND2X1 U632 ( .A(mem_28__3_), .B(n405), .Y(n409) );
  OAI211X1 U633 ( .C(n403), .D(n17), .A(n410), .B(n23), .Y(N782) );
  NAND2X1 U634 ( .A(mem_28__2_), .B(n405), .Y(n410) );
  OAI211X1 U635 ( .C(n403), .D(n25), .A(n411), .B(n31), .Y(N781) );
  NAND2X1 U636 ( .A(mem_28__1_), .B(n405), .Y(n411) );
  OAI211X1 U637 ( .C(n403), .D(n33), .A(n412), .B(n39), .Y(N780) );
  NAND2X1 U638 ( .A(mem_28__0_), .B(n405), .Y(n412) );
  NOR21XL U639 ( .B(n403), .A(n47), .Y(n405) );
  OAI22X1 U640 ( .A(n111), .B(n3), .C(n42), .D(n413), .Y(N779) );
  OAI21X1 U641 ( .B(gt_97_A_2_), .C(N693), .A(n342), .Y(n413) );
  NAND2X1 U642 ( .A(n365), .B(n402), .Y(n342) );
  OAI211X1 U643 ( .C(n414), .D(n50), .A(n415), .B(n56), .Y(N778) );
  NAND2X1 U644 ( .A(mem_29__7_), .B(n416), .Y(n415) );
  OAI211X1 U645 ( .C(n414), .D(n58), .A(n417), .B(n64), .Y(N777) );
  NAND2X1 U646 ( .A(mem_29__6_), .B(n416), .Y(n417) );
  OAI211X1 U647 ( .C(n414), .D(n66), .A(n418), .B(n72), .Y(N776) );
  NAND2X1 U648 ( .A(mem_29__5_), .B(n416), .Y(n418) );
  OAI211X1 U649 ( .C(n414), .D(n74), .A(n419), .B(n78), .Y(N775) );
  NAND2X1 U650 ( .A(mem_29__4_), .B(n416), .Y(n419) );
  OAI211X1 U651 ( .C(n414), .D(n9), .A(n420), .B(n15), .Y(N774) );
  NAND2X1 U652 ( .A(mem_29__3_), .B(n416), .Y(n420) );
  OAI211X1 U653 ( .C(n414), .D(n17), .A(n421), .B(n23), .Y(N773) );
  NAND2X1 U654 ( .A(mem_29__2_), .B(n416), .Y(n421) );
  OAI211X1 U655 ( .C(n414), .D(n25), .A(n422), .B(n31), .Y(N772) );
  NAND2X1 U656 ( .A(mem_29__1_), .B(n416), .Y(n422) );
  OAI211X1 U657 ( .C(n414), .D(n33), .A(n423), .B(n39), .Y(N771) );
  NAND2X1 U658 ( .A(mem_29__0_), .B(n416), .Y(n423) );
  NOR21XL U659 ( .B(n414), .A(n47), .Y(n416) );
  OAI22X1 U660 ( .A(n132), .B(n3), .C(n424), .D(n43), .Y(N770) );
  AOI21AX1 U661 ( .B(n134), .C(n378), .A(n425), .Y(n424) );
  OAI211X1 U662 ( .C(n426), .D(n50), .A(n427), .B(n56), .Y(N769) );
  NAND2X1 U663 ( .A(mem_30__7_), .B(n428), .Y(n427) );
  OAI211X1 U664 ( .C(n426), .D(n58), .A(n429), .B(n64), .Y(N768) );
  NAND2X1 U665 ( .A(mem_30__6_), .B(n428), .Y(n429) );
  OAI211X1 U666 ( .C(n426), .D(n66), .A(n430), .B(n72), .Y(N767) );
  NAND2X1 U667 ( .A(mem_30__5_), .B(n428), .Y(n430) );
  OAI211X1 U668 ( .C(n426), .D(n74), .A(n431), .B(n78), .Y(N766) );
  NAND2X1 U669 ( .A(mem_30__4_), .B(n428), .Y(n431) );
  OAI211X1 U670 ( .C(n426), .D(n9), .A(n432), .B(n15), .Y(N765) );
  NAND2X1 U671 ( .A(mem_30__3_), .B(n428), .Y(n432) );
  OAI211X1 U672 ( .C(n426), .D(n17), .A(n433), .B(n23), .Y(N764) );
  NAND2X1 U673 ( .A(mem_30__2_), .B(n428), .Y(n433) );
  OAI211X1 U674 ( .C(n426), .D(n25), .A(n434), .B(n31), .Y(N763) );
  NAND2X1 U675 ( .A(mem_30__1_), .B(n428), .Y(n434) );
  OAI211X1 U676 ( .C(n426), .D(n33), .A(n435), .B(n39), .Y(N762) );
  NAND2X1 U677 ( .A(mem_30__0_), .B(n428), .Y(n435) );
  NOR21XL U678 ( .B(n426), .A(n47), .Y(n428) );
  OAI22X1 U679 ( .A(n425), .B(n42), .C(n130), .D(n3), .Y(N761) );
  NAND2X1 U680 ( .A(n134), .B(n283), .Y(n130) );
  NOR2X1 U681 ( .A(n436), .B(n221), .Y(n134) );
  AOI21X1 U682 ( .B(n147), .C(n378), .A(N693), .Y(n425) );
  OAI211X1 U683 ( .C(n437), .D(n50), .A(n438), .B(n115), .Y(N760) );
  NAND2X1 U684 ( .A(mem_31__7_), .B(n439), .Y(n438) );
  OAI211X1 U685 ( .C(n437), .D(n58), .A(n440), .B(n119), .Y(N759) );
  NAND2X1 U686 ( .A(mem_31__6_), .B(n439), .Y(n440) );
  OAI211X1 U687 ( .C(n437), .D(n66), .A(n441), .B(n122), .Y(N758) );
  NAND2X1 U688 ( .A(mem_31__5_), .B(n439), .Y(n441) );
  OAI211X1 U689 ( .C(n437), .D(n74), .A(n442), .B(n78), .Y(N757) );
  NAND2X1 U690 ( .A(mem_31__4_), .B(n439), .Y(n442) );
  OAI211X1 U691 ( .C(n437), .D(n9), .A(n443), .B(n15), .Y(N756) );
  NAND2X1 U692 ( .A(mem_31__3_), .B(n439), .Y(n443) );
  OAI211X1 U693 ( .C(n437), .D(n17), .A(n444), .B(n23), .Y(N755) );
  NAND2X1 U694 ( .A(mem_31__2_), .B(n439), .Y(n444) );
  OAI211X1 U695 ( .C(n437), .D(n25), .A(n445), .B(n31), .Y(N754) );
  NAND2X1 U696 ( .A(mem_31__1_), .B(n439), .Y(n445) );
  OAI211X1 U697 ( .C(n437), .D(n33), .A(n446), .B(n39), .Y(N753) );
  NAND2X1 U698 ( .A(mem_31__0_), .B(n439), .Y(n446) );
  NOR21XL U699 ( .B(n437), .A(n47), .Y(n439) );
  ENOX1 U700 ( .A(n145), .B(n3), .C(n447), .D(n49), .Y(N752) );
  OAI21X1 U701 ( .B(n160), .C(n402), .A(n365), .Y(n447) );
  NAND2X1 U702 ( .A(n147), .B(n436), .Y(n145) );
  OAI211X1 U703 ( .C(n448), .D(n50), .A(n449), .B(n56), .Y(N751) );
  NAND2X1 U704 ( .A(mem_32__7_), .B(n450), .Y(n449) );
  OAI211X1 U705 ( .C(n448), .D(n58), .A(n451), .B(n64), .Y(N750) );
  NAND2X1 U706 ( .A(mem_32__6_), .B(n450), .Y(n451) );
  OAI211X1 U707 ( .C(n448), .D(n66), .A(n452), .B(n72), .Y(N749) );
  NAND2X1 U708 ( .A(mem_32__5_), .B(n450), .Y(n452) );
  OAI211X1 U709 ( .C(n448), .D(n74), .A(n453), .B(n78), .Y(N748) );
  NAND2X1 U710 ( .A(mem_32__4_), .B(n450), .Y(n453) );
  OAI211X1 U711 ( .C(n448), .D(n9), .A(n454), .B(n96), .Y(N747) );
  NAND2X1 U712 ( .A(mem_32__3_), .B(n450), .Y(n454) );
  OAI211X1 U713 ( .C(n448), .D(n17), .A(n455), .B(n100), .Y(N746) );
  NAND2X1 U714 ( .A(mem_32__2_), .B(n450), .Y(n455) );
  OAI211X1 U715 ( .C(n448), .D(n25), .A(n456), .B(n103), .Y(N745) );
  NAND2X1 U716 ( .A(mem_32__1_), .B(n450), .Y(n456) );
  OAI211X1 U717 ( .C(n448), .D(n33), .A(n457), .B(n39), .Y(N744) );
  NAND2X1 U718 ( .A(mem_32__0_), .B(n450), .Y(n457) );
  NOR21XL U719 ( .B(n448), .A(n47), .Y(n450) );
  OAI22X1 U720 ( .A(n42), .B(n365), .C(n160), .D(n376), .Y(N743) );
  INVX1 U721 ( .A(n402), .Y(n378) );
  NAND2X1 U722 ( .A(N1157), .B(N1159), .Y(n402) );
  NAND2X1 U723 ( .A(n147), .B(gt_97_A_0_), .Y(n160) );
  NOR2X1 U724 ( .A(n283), .B(n5), .Y(n147) );
  OAI211X1 U725 ( .C(n459), .D(n50), .A(n460), .B(n115), .Y(N742) );
  NAND2X1 U726 ( .A(mem_33__7_), .B(n461), .Y(n460) );
  OAI211X1 U727 ( .C(n459), .D(n58), .A(n462), .B(n119), .Y(N741) );
  NAND2X1 U728 ( .A(mem_33__6_), .B(n461), .Y(n462) );
  OAI211X1 U729 ( .C(n459), .D(n66), .A(n463), .B(n122), .Y(N740) );
  NAND2X1 U730 ( .A(mem_33__5_), .B(n461), .Y(n463) );
  OAI211X1 U731 ( .C(n459), .D(n74), .A(n464), .B(n78), .Y(N739) );
  NAND2X1 U732 ( .A(mem_33__4_), .B(n461), .Y(n464) );
  OAI211X1 U733 ( .C(n459), .D(n9), .A(n465), .B(n96), .Y(N738) );
  NAND2X1 U734 ( .A(mem_33__3_), .B(n461), .Y(n465) );
  OAI211X1 U735 ( .C(n459), .D(n17), .A(n466), .B(n100), .Y(N737) );
  NAND2X1 U736 ( .A(mem_33__2_), .B(n461), .Y(n466) );
  OAI211X1 U737 ( .C(n459), .D(n25), .A(n467), .B(n103), .Y(N736) );
  NAND2X1 U738 ( .A(mem_33__1_), .B(n461), .Y(n467) );
  OAI211X1 U739 ( .C(n459), .D(n33), .A(n468), .B(n39), .Y(N735) );
  NAND2X1 U740 ( .A(mem_33__0_), .B(n461), .Y(n468) );
  NOR21XL U741 ( .B(n459), .A(n47), .Y(n461) );
  OAI21BBX1 U742 ( .A(n49), .B(n469), .C(n458), .Y(N734) );
  NAND2X1 U743 ( .A(n471), .B(n472), .Y(n458) );
  AOI31X1 U744 ( .A(n472), .B(n257), .C(n318), .D(n365), .Y(n469) );
  INVX1 U745 ( .A(n172), .Y(n472) );
  OAI31XL U746 ( .A(n47), .B(add_101_B_0_), .C(n473), .D(n470), .Y(N733) );
  NAND21X1 U747 ( .B(n183), .A(n471), .Y(n470) );
  NOR43XL U748 ( .B(N693), .C(n269), .D(n318), .A(N1159), .Y(n471) );
  INVX1 U749 ( .A(full), .Y(add_101_B_0_) );
  INVX1 U750 ( .A(n365), .Y(N693) );
  AO22X1 U751 ( .A(N1040), .B(n474), .C(N1046), .D(n475), .Y(N1059) );
  AO22X1 U752 ( .A(N1039), .B(n474), .C(N1045), .D(n475), .Y(N1058) );
  AO22X1 U753 ( .A(N1038), .B(n474), .C(N1044), .D(n475), .Y(N1057) );
  AO22X1 U754 ( .A(N1037), .B(n474), .C(N1043), .D(n475), .Y(N1056) );
  AO22X1 U755 ( .A(N1036), .B(n474), .C(N1042), .D(n475), .Y(N1055) );
  AO22X1 U756 ( .A(N1035), .B(n474), .C(N1041), .D(n475), .Y(N1054) );
  NOR2X1 U757 ( .A(n476), .B(n477), .Y(n475) );
  NOR2X1 U758 ( .A(n477), .B(n478), .Y(n474) );
  NAND2X1 U759 ( .A(n477), .B(n479), .Y(N1053) );
  XNOR2XL U760 ( .A(n473), .B(n478), .Y(n477) );
  INVX1 U761 ( .A(n476), .Y(n478) );
  OAI211X1 U762 ( .C(n480), .D(n50), .A(n481), .B(n56), .Y(N1030) );
  NAND2X1 U763 ( .A(dat_7_1[7]), .B(n482), .Y(n481) );
  OAI211X1 U764 ( .C(n480), .D(n58), .A(n483), .B(n64), .Y(N1029) );
  NAND2X1 U765 ( .A(dat_7_1[6]), .B(n482), .Y(n483) );
  OAI211X1 U766 ( .C(n480), .D(n66), .A(n484), .B(n72), .Y(N1028) );
  NAND2X1 U767 ( .A(dat_7_1[5]), .B(n482), .Y(n484) );
  OAI211X1 U768 ( .C(n480), .D(n74), .A(n485), .B(n78), .Y(N1027) );
  NAND2X1 U769 ( .A(dat_7_1[4]), .B(n482), .Y(n485) );
  OAI211X1 U770 ( .C(n480), .D(n9), .A(n486), .B(n96), .Y(N1026) );
  NAND2X1 U771 ( .A(dat_7_1[3]), .B(n482), .Y(n486) );
  OAI211X1 U772 ( .C(n480), .D(n17), .A(n487), .B(n100), .Y(N1025) );
  NAND2X1 U773 ( .A(dat_7_1[2]), .B(n482), .Y(n487) );
  OAI211X1 U774 ( .C(n480), .D(n25), .A(n488), .B(n103), .Y(N1024) );
  NAND2X1 U775 ( .A(dat_7_1[1]), .B(n482), .Y(n488) );
  OAI211X1 U776 ( .C(n480), .D(n33), .A(n489), .B(n106), .Y(N1023) );
  NAND2X1 U777 ( .A(dat_7_1[0]), .B(n482), .Y(n489) );
  NOR21XL U778 ( .B(n480), .A(n47), .Y(n482) );
  OAI22X1 U779 ( .A(n490), .B(n42), .C(n1), .D(n172), .Y(N1022) );
  NAND3X1 U780 ( .A(n283), .B(n221), .C(n436), .Y(n172) );
  NOR2X1 U781 ( .A(n491), .B(gt_97_A_0_), .Y(n490) );
  OAI211X1 U782 ( .C(n492), .D(n50), .A(n493), .B(n56), .Y(N1021) );
  NAND2X1 U783 ( .A(dat_7_1[15]), .B(n494), .Y(n493) );
  OAI211X1 U784 ( .C(n492), .D(n58), .A(n495), .B(n64), .Y(N1020) );
  NAND2X1 U785 ( .A(dat_7_1[14]), .B(n494), .Y(n495) );
  OAI211X1 U786 ( .C(n492), .D(n66), .A(n496), .B(n72), .Y(N1019) );
  NAND2X1 U787 ( .A(dat_7_1[13]), .B(n494), .Y(n496) );
  OAI211X1 U788 ( .C(n492), .D(n74), .A(n497), .B(n78), .Y(N1018) );
  NAND2X1 U789 ( .A(dat_7_1[12]), .B(n494), .Y(n497) );
  OAI211X1 U790 ( .C(n492), .D(n9), .A(n498), .B(n13), .Y(N1017) );
  NAND2X1 U791 ( .A(dat_7_1[11]), .B(n494), .Y(n498) );
  OAI211X1 U792 ( .C(n492), .D(n17), .A(n499), .B(n21), .Y(N1016) );
  NAND2X1 U793 ( .A(dat_7_1[10]), .B(n494), .Y(n499) );
  OAI211X1 U794 ( .C(n492), .D(n25), .A(n500), .B(n29), .Y(N1015) );
  NAND2X1 U795 ( .A(dat_7_1[9]), .B(n494), .Y(n500) );
  OAI211X1 U796 ( .C(n492), .D(n33), .A(n501), .B(n106), .Y(N1014) );
  NAND2X1 U797 ( .A(dat_7_1[8]), .B(n494), .Y(n501) );
  NOR21XL U798 ( .B(n492), .A(n47), .Y(n494) );
  OAI22X1 U799 ( .A(n502), .B(n42), .C(n110), .D(n183), .Y(N1013) );
  INVX1 U800 ( .A(n491), .Y(n502) );
  NAND2X1 U801 ( .A(n108), .B(n283), .Y(n491) );
  OAI211X1 U802 ( .C(n503), .D(n50), .A(n504), .B(n56), .Y(N1012) );
  NAND2X1 U803 ( .A(dat_7_1[23]), .B(n505), .Y(n504) );
  OAI211X1 U804 ( .C(n503), .D(n58), .A(n506), .B(n64), .Y(N1011) );
  NAND2X1 U805 ( .A(dat_7_1[22]), .B(n505), .Y(n506) );
  OAI211X1 U806 ( .C(n503), .D(n66), .A(n507), .B(n72), .Y(N1010) );
  NAND2X1 U807 ( .A(dat_7_1[21]), .B(n505), .Y(n507) );
  OAI211X1 U808 ( .C(n503), .D(n74), .A(n508), .B(n78), .Y(N1009) );
  NAND2X1 U809 ( .A(dat_7_1[20]), .B(n505), .Y(n508) );
  OAI211X1 U810 ( .C(n503), .D(n9), .A(n13), .B(n509), .Y(N1008) );
  NAND2X1 U811 ( .A(dat_7_1[19]), .B(n505), .Y(n509) );
  NAND2X1 U812 ( .A(fifowdat[3]), .B(n41), .Y(n96) );
  MUX2IX1 U813 ( .D0(r_wdat[3]), .D1(prx_wdat[3]), .S(prx_psh), .Y(n95) );
  OAI211X1 U814 ( .C(n503), .D(n17), .A(n21), .B(n510), .Y(N1007) );
  NAND2X1 U815 ( .A(dat_7_1[18]), .B(n505), .Y(n510) );
  NAND2X1 U816 ( .A(fifowdat[2]), .B(n41), .Y(n100) );
  MUX2IX1 U817 ( .D0(r_wdat[2]), .D1(prx_wdat[2]), .S(prx_psh), .Y(n99) );
  OAI211X1 U818 ( .C(n503), .D(n25), .A(n29), .B(n511), .Y(N1006) );
  NAND2X1 U819 ( .A(dat_7_1[17]), .B(n505), .Y(n511) );
  NAND2X1 U820 ( .A(fifowdat[1]), .B(n41), .Y(n103) );
  MUX2IX1 U821 ( .D0(r_wdat[1]), .D1(prx_wdat[1]), .S(prx_psh), .Y(n102) );
  OAI211X1 U822 ( .C(n503), .D(n33), .A(n512), .B(n106), .Y(N1005) );
  NAND2X1 U823 ( .A(fifowdat[0]), .B(n41), .Y(n106) );
  NAND2X1 U824 ( .A(dat_7_1[16]), .B(n505), .Y(n512) );
  NOR21XL U825 ( .B(n503), .A(n47), .Y(n505) );
  MUX2IX1 U826 ( .D0(r_wdat[0]), .D1(prx_wdat[0]), .S(prx_psh), .Y(n105) );
  NAND2X1 U827 ( .A(n209), .B(n221), .Y(n111) );
  OAI22X1 U828 ( .A(n513), .B(n42), .C(n1), .D(n196), .Y(N1004) );
  NAND3X1 U829 ( .A(n436), .B(n221), .C(gt_97_A_1_), .Y(n196) );
  INVX1 U830 ( .A(n283), .Y(gt_97_A_1_) );
  NOR21XL U831 ( .B(n108), .A(n209), .Y(n513) );
  NOR2X1 U832 ( .A(n283), .B(n436), .Y(n209) );
  OAI211X1 U833 ( .C(n94), .D(n50), .A(n115), .B(n514), .Y(N1003) );
  NAND2X1 U834 ( .A(dat_7_1[31]), .B(n98), .Y(n514) );
  NAND2X1 U835 ( .A(fifowdat[7]), .B(n41), .Y(n115) );
  MUX2IX1 U836 ( .D0(r_wdat[7]), .D1(prx_wdat[7]), .S(prx_psh), .Y(n113) );
  OAI211X1 U837 ( .C(n94), .D(n58), .A(n119), .B(n515), .Y(N1002) );
  NAND2X1 U838 ( .A(dat_7_1[30]), .B(n98), .Y(n515) );
  NAND2X1 U839 ( .A(fifowdat[6]), .B(n41), .Y(n119) );
  OAI211X1 U840 ( .C(n94), .D(n66), .A(n122), .B(n516), .Y(N1001) );
  NAND2X1 U841 ( .A(dat_7_1[29]), .B(n98), .Y(n516) );
  NAND2X1 U842 ( .A(fifowdat[5]), .B(n41), .Y(n122) );
  MUX2IX1 U843 ( .D0(r_wdat[5]), .D1(prx_wdat[5]), .S(prx_psh), .Y(n120) );
  OAI211X1 U844 ( .C(n94), .D(n74), .A(n517), .B(n78), .Y(N1000) );
  NAND2X1 U845 ( .A(fifowdat[4]), .B(n41), .Y(n125) );
  NAND2X1 U846 ( .A(dat_7_1[28]), .B(n98), .Y(n517) );
  NOR21XL U847 ( .B(n94), .A(n44), .Y(n98) );
  OAI21X1 U848 ( .B(n90), .C(n518), .A(n519), .Y(n476) );
  NOR2X1 U849 ( .A(n146), .B(gt_97_A_2_), .Y(n108) );
  NAND3X1 U850 ( .A(n436), .B(n283), .C(gt_97_A_2_), .Y(n132) );
  INVX1 U851 ( .A(n221), .Y(gt_97_A_2_) );
  INVX1 U852 ( .A(n146), .Y(n159) );
  NAND2X1 U853 ( .A(n222), .B(n257), .Y(n146) );
  INVX1 U854 ( .A(n245), .Y(n222) );
  NAND2X1 U855 ( .A(n318), .B(n365), .Y(n245) );
  NOR2X1 U856 ( .A(n473), .B(full), .Y(n269) );
  INVX1 U857 ( .A(fifopsh), .Y(n473) );
  OAI21X1 U858 ( .B(n90), .C(n520), .A(n521), .Y(fifopsh) );
  NOR2X1 U859 ( .A(r_unlock), .B(ps_locked), .Y(n90) );
  NOR43XL U860 ( .B(n519), .C(n479), .D(n521), .A(n522), .Y(ps_locked) );
  AOI21X1 U861 ( .B(i_lockena), .C(n92), .A(locked), .Y(n522) );
  NAND2X1 U862 ( .A(n520), .B(n518), .Y(n92) );
  INVX1 U863 ( .A(r_pop), .Y(n518) );
  INVX1 U864 ( .A(r_psh), .Y(n520) );
  INVX1 U865 ( .A(prx_psh), .Y(n521) );
  NOR21XL U866 ( .B(srstz), .A(r_fiforst), .Y(n479) );
  INVX1 U867 ( .A(ptx_pop), .Y(n519) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_1 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_2 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_3 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_4 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_5 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_6 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_7 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_8 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_9 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_10 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_11 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_12 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_13 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_14 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_15 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_16 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_17 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_18 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_19 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_20 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_21 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_22 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_23 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_24 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_25 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_26 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_27 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_28 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_29 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_30 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_31 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_32 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_33 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_34 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyff_DEPTH_NUM34_DEPTH_NBT6_0 ( CLK, EN, ENCLK, 
        TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module phycrc_a0 ( crc32_3_0, rx_good, i_shfidat, i_start, i_shfi4, i_shfo4, 
        clk );
  output [3:0] crc32_3_0;
  input [3:0] i_shfidat;
  input i_start, i_shfi4, i_shfo4, clk;
  output rx_good;
  wire   N188, N189, N190, N191, N192, N193, N194, N195, N196, N197, N198,
         N199, N200, N201, N202, N203, N204, N205, N206, N207, N208, N209,
         N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220,
         net10566, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n1, n2, n3, n4, n5, n6, n7, n8,
         n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n55, n119, n120,
         n121, n122, n124, n125, n126, n127;
  wire   [31:0] crc32_r;

  SNPS_CLOCK_GATE_HIGH_phycrc_a0 clk_gate_crc32_r_reg ( .CLK(clk), .EN(N188), 
        .ENCLK(net10566), .TE(1'b0) );
  DFFQX1 crc32_r_reg_26_ ( .D(N215), .C(net10566), .Q(crc32_r[26]) );
  DFFQX1 crc32_r_reg_16_ ( .D(N205), .C(net10566), .Q(crc32_r[16]) );
  DFFQX1 crc32_r_reg_4_ ( .D(N193), .C(net10566), .Q(crc32_r[4]) );
  DFFQX1 crc32_r_reg_3_ ( .D(N192), .C(net10566), .Q(crc32_r[3]) );
  DFFQX1 crc32_r_reg_25_ ( .D(N214), .C(net10566), .Q(crc32_r[25]) );
  DFFQX1 crc32_r_reg_24_ ( .D(N213), .C(net10566), .Q(crc32_r[24]) );
  DFFQX1 crc32_r_reg_27_ ( .D(N216), .C(net10566), .Q(crc32_r[27]) );
  DFFQX1 crc32_r_reg_17_ ( .D(N206), .C(net10566), .Q(crc32_r[17]) );
  DFFQX1 crc32_r_reg_11_ ( .D(N200), .C(net10566), .Q(crc32_r[11]) );
  DFFQX1 crc32_r_reg_15_ ( .D(N204), .C(net10566), .Q(crc32_r[15]) );
  DFFQX1 crc32_r_reg_0_ ( .D(N189), .C(net10566), .Q(crc32_r[0]) );
  DFFQX1 crc32_r_reg_8_ ( .D(N197), .C(net10566), .Q(crc32_r[8]) );
  DFFQX1 crc32_r_reg_5_ ( .D(N194), .C(net10566), .Q(crc32_r[5]) );
  DFFQX1 crc32_r_reg_1_ ( .D(N190), .C(net10566), .Q(crc32_r[1]) );
  DFFQX1 crc32_r_reg_10_ ( .D(N199), .C(net10566), .Q(crc32_r[10]) );
  DFFQX1 crc32_r_reg_6_ ( .D(N195), .C(net10566), .Q(crc32_r[6]) );
  DFFQX1 crc32_r_reg_12_ ( .D(N201), .C(net10566), .Q(crc32_r[12]) );
  DFFQX1 crc32_r_reg_14_ ( .D(N203), .C(net10566), .Q(crc32_r[14]) );
  DFFQX1 crc32_r_reg_18_ ( .D(N207), .C(net10566), .Q(crc32_r[18]) );
  DFFQX1 crc32_r_reg_9_ ( .D(N198), .C(net10566), .Q(crc32_r[9]) );
  DFFQX1 crc32_r_reg_21_ ( .D(N210), .C(net10566), .Q(crc32_r[21]) );
  DFFQX1 crc32_r_reg_20_ ( .D(N209), .C(net10566), .Q(crc32_r[20]) );
  DFFQX1 crc32_r_reg_7_ ( .D(N196), .C(net10566), .Q(crc32_r[7]) );
  DFFQX1 crc32_r_reg_22_ ( .D(N211), .C(net10566), .Q(crc32_r[22]) );
  DFFQX1 crc32_r_reg_13_ ( .D(N202), .C(net10566), .Q(crc32_r[13]) );
  DFFQX1 crc32_r_reg_2_ ( .D(N191), .C(net10566), .Q(crc32_r[2]) );
  DFFQX1 crc32_r_reg_23_ ( .D(N212), .C(net10566), .Q(crc32_r[23]) );
  DFFQX1 crc32_r_reg_28_ ( .D(N217), .C(net10566), .Q(crc32_r[28]) );
  DFFQX1 crc32_r_reg_29_ ( .D(N218), .C(net10566), .Q(crc32_r[29]) );
  DFFQX1 crc32_r_reg_19_ ( .D(N208), .C(net10566), .Q(crc32_r[19]) );
  DFFQX1 crc32_r_reg_31_ ( .D(N220), .C(net10566), .Q(crc32_r[31]) );
  DFFQX1 crc32_r_reg_30_ ( .D(N219), .C(net10566), .Q(crc32_r[30]) );
  BUFX3 U3 ( .A(n59), .Y(n1) );
  NOR2X1 U4 ( .A(n13), .B(n78), .Y(n2) );
  INVX1 U5 ( .A(n13), .Y(n3) );
  INVX1 U6 ( .A(n78), .Y(n4) );
  INVX1 U7 ( .A(n14), .Y(n5) );
  XNOR2XL U8 ( .A(i_shfidat[3]), .B(n117), .Y(n69) );
  INVX1 U9 ( .A(n75), .Y(n6) );
  XNOR2XL U10 ( .A(i_shfidat[1]), .B(n114), .Y(n48) );
  XNOR2XL U11 ( .A(i_shfidat[2]), .B(n116), .Y(n53) );
  NAND2X1 U12 ( .A(n9), .B(n57), .Y(N188) );
  NAND21X1 U13 ( .B(n9), .A(n1), .Y(n43) );
  INVX1 U14 ( .A(n75), .Y(n12) );
  NAND2X1 U15 ( .A(i_shfo4), .B(n11), .Y(n8) );
  NAND2X1 U16 ( .A(i_shfo4), .B(n9), .Y(n57) );
  INVX1 U17 ( .A(n7), .Y(n9) );
  INVX1 U18 ( .A(n7), .Y(n11) );
  INVX1 U19 ( .A(n7), .Y(n10) );
  NOR2X1 U20 ( .A(n17), .B(i_start), .Y(n59) );
  NOR2X1 U21 ( .A(n16), .B(i_start), .Y(n65) );
  INVX1 U22 ( .A(i_start), .Y(n13) );
  NOR2X1 U23 ( .A(i_shfi4), .B(n9), .Y(n75) );
  AOI21X1 U24 ( .B(n15), .C(n3), .A(n75), .Y(n52) );
  AOI21X1 U25 ( .B(n14), .C(n3), .A(n75), .Y(n72) );
  NOR2X1 U26 ( .A(n9), .B(i_start), .Y(n49) );
  NOR2X1 U27 ( .A(n75), .B(n66), .Y(n47) );
  OAI21X1 U28 ( .B(n11), .C(n14), .A(n6), .Y(N189) );
  OAI21X1 U29 ( .B(n11), .C(n112), .A(n6), .Y(N191) );
  XNOR2XL U30 ( .A(n14), .B(n113), .Y(n112) );
  XNOR2XL U31 ( .A(n15), .B(n16), .Y(n113) );
  OAI21X1 U32 ( .B(n11), .C(n109), .A(n6), .Y(N192) );
  XNOR2XL U33 ( .A(n15), .B(n110), .Y(n109) );
  XNOR2XL U34 ( .A(n16), .B(n4), .Y(n110) );
  OAI21X1 U35 ( .B(n11), .C(n115), .A(n6), .Y(N190) );
  XNOR2XL U36 ( .A(n14), .B(n15), .Y(n115) );
  OR2X1 U37 ( .A(i_start), .B(i_shfi4), .Y(n7) );
  NOR2X1 U38 ( .A(n75), .B(n60), .Y(n45) );
  INVX1 U39 ( .A(n48), .Y(n16) );
  INVX1 U40 ( .A(n78), .Y(n17) );
  NOR2X1 U41 ( .A(n13), .B(n78), .Y(n60) );
  NOR2X1 U42 ( .A(n13), .B(n48), .Y(n66) );
  OA21X1 U43 ( .B(n11), .C(n78), .A(n57), .Y(n44) );
  INVX1 U44 ( .A(n53), .Y(n15) );
  INVX1 U45 ( .A(n69), .Y(n14) );
  OAI21X1 U46 ( .B(n11), .C(n53), .A(n57), .Y(n54) );
  OAI21X1 U47 ( .B(n11), .C(n48), .A(n57), .Y(n50) );
  OAI21X1 U48 ( .B(n11), .C(n69), .A(n8), .Y(n73) );
  NOR4XL U49 ( .A(n18), .B(n119), .C(n30), .D(n21), .Y(n38) );
  NOR4XL U50 ( .A(n120), .B(n31), .C(n121), .D(n29), .Y(n37) );
  NOR4XL U51 ( .A(n19), .B(n24), .C(n126), .D(n20), .Y(n35) );
  NOR2X1 U52 ( .A(crc32_r[30]), .B(i_start), .Y(n114) );
  XNOR2XL U53 ( .A(i_shfidat[0]), .B(n111), .Y(n78) );
  NOR2X1 U54 ( .A(crc32_r[31]), .B(i_start), .Y(n111) );
  OAI221X1 U55 ( .A(n10), .B(n87), .C(n57), .D(n127), .E(n12), .Y(N200) );
  XNOR2XL U56 ( .A(n88), .B(n69), .Y(n87) );
  XNOR2XL U57 ( .A(n89), .B(n53), .Y(n88) );
  AOI221XL U58 ( .A(crc32_r[7]), .B(n17), .C(n59), .D(n127), .E(n60), .Y(n89)
         );
  OAI221X1 U59 ( .A(n10), .B(n103), .C(n29), .D(n8), .E(n12), .Y(N194) );
  XNOR2XL U60 ( .A(n104), .B(n69), .Y(n103) );
  XNOR2XL U61 ( .A(n105), .B(n53), .Y(n104) );
  AOI221XL U62 ( .A(crc32_r[1]), .B(n17), .C(n59), .D(n29), .E(n2), .Y(n105)
         );
  OAI221X1 U63 ( .A(n10), .B(n84), .C(n20), .D(n8), .E(n12), .Y(N201) );
  XNOR2XL U64 ( .A(n85), .B(n69), .Y(n84) );
  XNOR2XL U65 ( .A(n86), .B(n53), .Y(n85) );
  AOI221XL U66 ( .A(crc32_r[8]), .B(n16), .C(n65), .D(n20), .E(n66), .Y(n86)
         );
  OAI221X1 U67 ( .A(n10), .B(n95), .C(n19), .D(n57), .E(n12), .Y(N197) );
  XNOR2XL U68 ( .A(n96), .B(n69), .Y(n95) );
  XNOR2XL U69 ( .A(n97), .B(n53), .Y(n96) );
  AOI221XL U70 ( .A(crc32_r[4]), .B(n17), .C(n59), .D(n19), .E(n60), .Y(n97)
         );
  OAI221X1 U71 ( .A(n10), .B(n98), .C(n124), .D(n8), .E(n12), .Y(N196) );
  XNOR2XL U72 ( .A(n99), .B(n69), .Y(n98) );
  XNOR2XL U73 ( .A(n100), .B(n48), .Y(n99) );
  AOI221XL U74 ( .A(crc32_r[3]), .B(n17), .C(n59), .D(n124), .E(n60), .Y(n100)
         );
  OAI221X1 U75 ( .A(n10), .B(n90), .C(n126), .D(n57), .E(n12), .Y(N199) );
  XNOR2XL U76 ( .A(n91), .B(n69), .Y(n90) );
  XNOR2XL U77 ( .A(n92), .B(n48), .Y(n91) );
  AOI221XL U78 ( .A(crc32_r[6]), .B(n17), .C(n59), .D(n126), .E(n2), .Y(n92)
         );
  OAI221X1 U79 ( .A(n10), .B(n106), .C(n18), .D(n8), .E(n12), .Y(N193) );
  XNOR2XL U80 ( .A(n107), .B(n69), .Y(n106) );
  XNOR2XL U81 ( .A(n108), .B(n48), .Y(n107) );
  AOI221XL U82 ( .A(crc32_r[0]), .B(n17), .C(n59), .D(n18), .E(n60), .Y(n108)
         );
  OAI221X1 U83 ( .A(n9), .B(n81), .C(n8), .D(n25), .E(n12), .Y(N202) );
  XNOR2XL U84 ( .A(n82), .B(n53), .Y(n81) );
  XNOR2XL U85 ( .A(n83), .B(n48), .Y(n82) );
  AOI221XL U86 ( .A(crc32_r[9]), .B(n17), .C(n59), .D(n25), .E(n2), .Y(n83) );
  OAI221X1 U87 ( .A(n9), .B(n67), .C(n57), .D(n32), .E(n12), .Y(N212) );
  INVX1 U88 ( .A(crc32_r[19]), .Y(n32) );
  XNOR2XL U89 ( .A(n68), .B(n69), .Y(n67) );
  XNOR2XL U90 ( .A(n70), .B(n53), .Y(n68) );
  OAI221X1 U91 ( .A(n10), .B(n56), .C(n122), .D(n8), .E(n12), .Y(N215) );
  XNOR2XL U92 ( .A(n58), .B(n14), .Y(n56) );
  AOI221XL U93 ( .A(crc32_r[22]), .B(n4), .C(n1), .D(n122), .E(n2), .Y(n58) );
  INVX1 U94 ( .A(crc32_r[22]), .Y(n122) );
  OAI221X1 U95 ( .A(n9), .B(n79), .C(n119), .D(n57), .E(n6), .Y(N203) );
  XNOR2XL U96 ( .A(n80), .B(n16), .Y(n79) );
  AOI221XL U97 ( .A(crc32_r[10]), .B(n17), .C(n59), .D(n119), .E(n2), .Y(n80)
         );
  OAI221X1 U98 ( .A(n10), .B(n93), .C(n24), .D(n8), .E(n6), .Y(N198) );
  XNOR2XL U99 ( .A(n94), .B(n15), .Y(n93) );
  AOI221XL U100 ( .A(crc32_r[5]), .B(n16), .C(n65), .D(n24), .E(n66), .Y(n94)
         );
  OAI221X1 U101 ( .A(n10), .B(n101), .C(n8), .D(n125), .E(n6), .Y(N195) );
  XNOR2XL U102 ( .A(n102), .B(n15), .Y(n101) );
  AOI221XL U103 ( .A(crc32_r[2]), .B(n16), .C(n65), .D(n125), .E(n66), .Y(n102) );
  INVX1 U104 ( .A(crc32_r[2]), .Y(n125) );
  OAI221X1 U105 ( .A(n9), .B(n61), .C(n57), .D(n27), .E(n6), .Y(N214) );
  XNOR2XL U106 ( .A(n62), .B(n16), .Y(n61) );
  AOI221XL U107 ( .A(crc32_r[21]), .B(n17), .C(n59), .D(n27), .E(n60), .Y(n62)
         );
  INVX1 U108 ( .A(crc32_r[21]), .Y(n27) );
  OAI221X1 U109 ( .A(n9), .B(n63), .C(n8), .D(n22), .E(n6), .Y(N213) );
  XNOR2XL U110 ( .A(n64), .B(n15), .Y(n63) );
  AOI221XL U111 ( .A(crc32_r[20]), .B(n16), .C(n65), .D(n22), .E(n66), .Y(n64)
         );
  INVX1 U112 ( .A(crc32_r[20]), .Y(n22) );
  NOR2X1 U113 ( .A(crc32_r[29]), .B(i_start), .Y(n116) );
  NOR2X1 U114 ( .A(crc32_r[28]), .B(i_start), .Y(n117) );
  NAND2X1 U115 ( .A(n71), .B(n72), .Y(N211) );
  AOI32X1 U116 ( .A(n49), .B(n121), .C(n5), .D(crc32_r[18]), .E(n73), .Y(n71)
         );
  NAND2X1 U117 ( .A(n74), .B(n47), .Y(N207) );
  AOI32X1 U118 ( .A(n48), .B(n120), .C(n49), .D(crc32_r[14]), .E(n50), .Y(n74)
         );
  NAND2X1 U119 ( .A(n51), .B(n52), .Y(N216) );
  AOI32X1 U120 ( .A(n49), .B(n55), .C(n53), .D(crc32_r[23]), .E(n54), .Y(n51)
         );
  INVX1 U121 ( .A(crc32_r[23]), .Y(n55) );
  NAND2X1 U122 ( .A(n76), .B(n52), .Y(N206) );
  AOI32X1 U123 ( .A(n49), .B(n26), .C(n53), .D(crc32_r[13]), .E(n54), .Y(n76)
         );
  INVX1 U124 ( .A(crc32_r[13]), .Y(n26) );
  NAND2X1 U125 ( .A(n46), .B(n47), .Y(N217) );
  AOI32X1 U126 ( .A(n48), .B(n23), .C(n49), .D(crc32_r[24]), .E(n50), .Y(n46)
         );
  INVX1 U127 ( .A(crc32_r[24]), .Y(n23) );
  NAND2X1 U128 ( .A(n77), .B(n72), .Y(N205) );
  AOI32X1 U129 ( .A(n49), .B(n21), .C(n5), .D(crc32_r[12]), .E(n73), .Y(n77)
         );
  OAI221X1 U130 ( .A(crc32_r[15]), .B(n43), .C(n44), .D(n31), .E(n45), .Y(N208) );
  OAI221X1 U131 ( .A(crc32_r[11]), .B(n43), .C(n44), .D(n30), .E(n45), .Y(N204) );
  OAI221X1 U132 ( .A(crc32_r[25]), .B(n43), .C(n44), .D(n28), .E(n45), .Y(N218) );
  INVX1 U133 ( .A(crc32_r[25]), .Y(n28) );
  NOR2X1 U134 ( .A(crc32_r[19]), .B(i_start), .Y(n70) );
  OAI21BBX1 U135 ( .A(N188), .B(crc32_r[26]), .C(n13), .Y(N219) );
  OAI21BBX1 U136 ( .A(N188), .B(crc32_r[27]), .C(n13), .Y(N220) );
  OAI21BBX1 U137 ( .A(N188), .B(crc32_r[17]), .C(n13), .Y(N210) );
  OAI21BBX1 U138 ( .A(N188), .B(crc32_r[16]), .C(n13), .Y(N209) );
  NOR2X1 U139 ( .A(n33), .B(n34), .Y(rx_good) );
  NAND4X1 U140 ( .A(n35), .B(n36), .C(n37), .D(n38), .Y(n34) );
  NAND4X1 U141 ( .A(n39), .B(n40), .C(n41), .D(n42), .Y(n33) );
  NOR43XL U142 ( .B(crc32_r[24]), .C(crc32_r[25]), .D(crc32_r[26]), .A(n124), 
        .Y(n36) );
  NOR4XL U143 ( .A(crc32_r[9]), .B(crc32_r[7]), .C(crc32_r[2]), .D(crc32_r[29]), .Y(n42) );
  NOR4XL U144 ( .A(crc32_r[28]), .B(crc32_r[27]), .C(crc32_r[23]), .D(
        crc32_r[22]), .Y(n41) );
  NOR4XL U145 ( .A(crc32_r[21]), .B(crc32_r[20]), .C(crc32_r[19]), .D(
        crc32_r[17]), .Y(n40) );
  NOR4XL U146 ( .A(crc32_r[16]), .B(crc32_r[13]), .C(crc32_3_0[1]), .D(
        crc32_3_0[0]), .Y(n39) );
  INVX1 U147 ( .A(crc32_r[30]), .Y(crc32_3_0[1]) );
  INVX1 U148 ( .A(crc32_r[31]), .Y(crc32_3_0[0]) );
  INVX1 U149 ( .A(crc32_r[6]), .Y(n126) );
  INVX1 U150 ( .A(crc32_r[1]), .Y(n29) );
  INVX1 U151 ( .A(crc32_r[8]), .Y(n20) );
  INVX1 U152 ( .A(crc32_r[10]), .Y(n119) );
  INVX1 U153 ( .A(crc32_r[5]), .Y(n24) );
  INVX1 U154 ( .A(crc32_r[0]), .Y(n18) );
  INVX1 U155 ( .A(crc32_r[18]), .Y(n121) );
  INVX1 U156 ( .A(crc32_r[12]), .Y(n21) );
  INVX1 U157 ( .A(crc32_r[14]), .Y(n120) );
  INVX1 U158 ( .A(crc32_r[11]), .Y(n30) );
  INVX1 U159 ( .A(crc32_r[15]), .Y(n31) );
  INVX1 U160 ( .A(crc32_r[28]), .Y(crc32_3_0[3]) );
  INVX1 U161 ( .A(crc32_r[29]), .Y(crc32_3_0[2]) );
  INVX1 U162 ( .A(crc32_r[3]), .Y(n124) );
  INVX1 U163 ( .A(crc32_r[4]), .Y(n19) );
  INVX1 U164 ( .A(crc32_r[7]), .Y(n127) );
  INVX1 U165 ( .A(crc32_r[9]), .Y(n25) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phycrc_a0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module phytx_a0 ( r_txnumk, r_txendk, r_txshrt, r_txauto, prx_cccnt, ptx_txact, 
        ptx_cc, ptx_goidle, ptx_fifopop, ptx_pspyld, i_rdat, i_txreq, i_one, 
        ptx_crcstart, ptx_crcshfi4, ptx_crcshfo4, ptx_crcsidat, ptx_fsm, 
        pcc_crc30, clk, srstz );
  input [4:0] r_txnumk;
  input [6:0] r_txauto;
  input [1:0] prx_cccnt;
  input [7:0] i_rdat;
  output [3:0] ptx_crcsidat;
  output [2:0] ptx_fsm;
  input [3:0] pcc_crc30;
  input r_txendk, r_txshrt, i_txreq, i_one, clk, srstz;
  output ptx_txact, ptx_cc, ptx_goidle, ptx_fifopop, ptx_pspyld, ptx_crcstart,
         ptx_crcshfi4, ptx_crcshfo4;
  wire   N45, hinib, N251, N252, N253, N254, N255, N264, N265, N266, N267,
         N268, N269, N270, N271, N272, N273, N297, N298, N299, net10588,
         net10594, n237, n238, n1, n2, n3, n4, n5, n6, n7, n8, n9, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250;
  wire   [4:0] bytcnt;
  wire   [3:0] bitcnt;
  wire   [3:0] encout;
  wire   [4:2] add_104_carry;

  SNPS_CLOCK_GATE_HIGH_phytx_a0_0 clk_gate_bitcnt_reg ( .CLK(clk), .EN(N251), 
        .ENCLK(net10588), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_phytx_a0_1 clk_gate_bytcnt_reg ( .CLK(clk), .EN(N268), 
        .ENCLK(net10594), .TE(1'b0) );
  DFFQX1 ptx_cc_reg ( .D(n238), .C(clk), .Q(ptx_cc) );
  DFFQX1 bitcnt_reg_3_ ( .D(N255), .C(net10588), .Q(bitcnt[3]) );
  DFFQX1 bitcnt_reg_0_ ( .D(N252), .C(net10588), .Q(bitcnt[0]) );
  DFFQX1 bitcnt_reg_1_ ( .D(N253), .C(net10588), .Q(bitcnt[1]) );
  DFFQX1 bitcnt_reg_2_ ( .D(N254), .C(net10588), .Q(bitcnt[2]) );
  DFFQX1 cs_txph_reg_2_ ( .D(N299), .C(clk), .Q(ptx_fsm[2]) );
  DFFQX1 cs_txph_reg_1_ ( .D(N298), .C(clk), .Q(ptx_fsm[1]) );
  DFFQX1 cs_txph_reg_0_ ( .D(N297), .C(clk), .Q(ptx_fsm[0]) );
  DFFQX1 bytcnt_reg_4_ ( .D(N273), .C(net10594), .Q(bytcnt[4]) );
  DFFQX1 bytcnt_reg_2_ ( .D(N271), .C(net10594), .Q(bytcnt[2]) );
  DFFQX1 bytcnt_reg_3_ ( .D(N272), .C(net10594), .Q(bytcnt[3]) );
  DFFQX1 bytcnt_reg_1_ ( .D(N270), .C(net10594), .Q(bytcnt[1]) );
  HAD1XL add_104_U1_1_2 ( .A(bytcnt[2]), .B(add_104_carry[2]), .CO(
        add_104_carry[3]), .SO(N265) );
  HAD1XL add_104_U1_1_1 ( .A(bytcnt[1]), .B(bytcnt[0]), .CO(add_104_carry[2]), 
        .SO(N264) );
  HAD1XL add_104_U1_1_3 ( .A(bytcnt[3]), .B(add_104_carry[3]), .CO(
        add_104_carry[4]), .SO(N266) );
  DFFQX1 bytcnt_reg_0_ ( .D(N269), .C(net10594), .Q(bytcnt[0]) );
  DFFQX1 hinib_reg ( .D(n237), .C(net10588), .Q(hinib) );
  NOR4X2 U3 ( .A(n132), .B(n131), .C(n190), .D(n6), .Y(n5) );
  XOR2X2 U4 ( .A(n130), .B(bitcnt[1]), .Y(n131) );
  INVX1 U5 ( .A(i_rdat[7]), .Y(n124) );
  INVX1 U6 ( .A(i_rdat[0]), .Y(n150) );
  INVX1 U7 ( .A(i_rdat[4]), .Y(n128) );
  AO21X1 U8 ( .B(n29), .C(n148), .A(n217), .Y(n215) );
  NAND5XL U9 ( .A(n204), .B(bytcnt[0]), .C(n136), .D(n135), .E(n134), .Y(n147)
         );
  NAND6XL U10 ( .A(n154), .B(n153), .C(n152), .D(n151), .E(n150), .F(n149), 
        .Y(n221) );
  NOR6XL U11 ( .A(i_rdat[5]), .B(bytcnt[1]), .C(i_rdat[4]), .D(n148), .E(n155), 
        .F(n147), .Y(n149) );
  INVX1 U12 ( .A(i_rdat[6]), .Y(n19) );
  INVX1 U13 ( .A(n43), .Y(n1) );
  MUX2X1 U14 ( .D0(n152), .D1(n124), .S(hinib), .Y(n52) );
  MUX2X1 U15 ( .D0(n150), .D1(n128), .S(hinib), .Y(n32) );
  MUX2IX1 U16 ( .D0(n153), .D1(n19), .S(hinib), .Y(ptx_crcsidat[2]) );
  INVX1 U17 ( .A(n52), .Y(ptx_crcsidat[3]) );
  NAND21X1 U18 ( .B(r_txnumk[1]), .A(bytcnt[1]), .Y(n207) );
  NOR2X1 U19 ( .A(n197), .B(n217), .Y(n2) );
  INVX1 U20 ( .A(bitcnt[3]), .Y(n6) );
  AOI22BXL U21 ( .B(bytcnt[3]), .A(r_txnumk[3]), .D(bytcnt[2]), .C(r_txnumk[2]), .Y(n22) );
  NAND42XL U22 ( .C(bitcnt[3]), .D(n131), .A(n4), .B(bitcnt[2]), .Y(n129) );
  NAND21XL U23 ( .B(n204), .A(n203), .Y(n206) );
  NAND21XL U24 ( .B(n145), .A(n130), .Y(n31) );
  GEN2X1 U25 ( .D(n36), .E(n30), .C(n126), .B(n77), .A(n145), .Y(n130) );
  MUX2BX1 U26 ( .D0(ptx_crcsidat[3]), .D1(n21), .S(ptx_crcsidat[2]), .Y(n30)
         );
  OAI31XL U27 ( .A(n133), .B(n215), .C(n203), .D(n143), .Y(n185) );
  AOI31XL U28 ( .A(n128), .B(n127), .C(n151), .D(n126), .Y(n133) );
  INVXL U29 ( .A(i_rdat[1]), .Y(n154) );
  INVXL U30 ( .A(r_txauto[6]), .Y(n126) );
  OA21XL U31 ( .B(r_txnumk[0]), .C(n223), .A(n207), .Y(n213) );
  AND4XL U32 ( .A(n211), .B(n210), .C(n209), .D(n208), .Y(n212) );
  NAND32XL U33 ( .B(n139), .C(n217), .A(n185), .Y(n173) );
  NAND21XL U34 ( .B(r_txauto[6]), .A(n37), .Y(n103) );
  NAND32XL U35 ( .B(n32), .C(n126), .A(n37), .Y(n65) );
  AO21XL U36 ( .B(i_rdat[1]), .C(n112), .A(n49), .Y(n56) );
  OR4X1 U37 ( .A(n161), .B(n105), .C(n41), .D(n3), .Y(encout[0]) );
  AOI21X1 U38 ( .B(n241), .C(n40), .A(n155), .Y(n3) );
  OAI221XL U39 ( .A(n104), .B(n155), .C(n103), .D(n128), .E(n102), .Y(n107) );
  NAND3XL U40 ( .A(r_txauto[6]), .B(n52), .C(n130), .Y(n9) );
  INVXL U41 ( .A(n32), .Y(ptx_crcsidat[0]) );
  XNOR2XL U42 ( .A(n130), .B(bitcnt[0]), .Y(n4) );
  NAND21XL U43 ( .B(r_txnumk[2]), .A(bytcnt[2]), .Y(n214) );
  OAI211XL U44 ( .C(n2), .D(n183), .A(n11), .B(n182), .Y(n243) );
  MUX2XL U45 ( .D0(n201), .D1(n1), .S(n200), .Y(n237) );
  AND3XL U46 ( .A(n227), .B(n211), .C(n197), .Y(n201) );
  INVXL U47 ( .A(n36), .Y(ptx_crcsidat[1]) );
  INVXL U48 ( .A(bytcnt[1]), .Y(n138) );
  MUX2BXL U49 ( .D0(bitcnt[1]), .D1(n7), .S(n1), .Y(N45) );
  XNOR2XL U50 ( .A(n131), .B(n88), .Y(n7) );
  OAI221XL U51 ( .A(hinib), .B(n45), .C(n232), .D(n44), .E(n236), .Y(n46) );
  MUX2XL U52 ( .D0(bytcnt[0]), .D1(hinib), .S(r_txauto[0]), .Y(n71) );
  OA22XL U53 ( .A(n229), .B(n230), .C(bytcnt[0]), .D(n228), .Y(n72) );
  OAI211XL U54 ( .C(bytcnt[0]), .D(hinib), .A(n240), .B(n20), .Y(n73) );
  MUX2XL U55 ( .D0(n68), .D1(n67), .S(hinib), .Y(n69) );
  INVXL U56 ( .A(bytcnt[0]), .Y(n223) );
  INVXL U57 ( .A(hinib), .Y(n43) );
  NAND2XL U58 ( .A(bytcnt[0]), .B(hinib), .Y(n240) );
  NAND21X1 U59 ( .B(n193), .A(n191), .Y(N251) );
  INVX1 U60 ( .A(n99), .Y(n38) );
  INVX1 U61 ( .A(n51), .Y(n82) );
  INVX1 U62 ( .A(n42), .Y(n95) );
  INVX1 U63 ( .A(n62), .Y(n54) );
  INVX1 U64 ( .A(srstz), .Y(n18) );
  INVX1 U65 ( .A(n143), .Y(n204) );
  INVX1 U66 ( .A(n185), .Y(n197) );
  INVX1 U67 ( .A(n188), .Y(n193) );
  NAND21X1 U68 ( .B(n187), .A(n191), .Y(n188) );
  INVX1 U69 ( .A(n186), .Y(n191) );
  NAND32X1 U70 ( .B(i_txreq), .C(n185), .A(n184), .Y(n186) );
  INVX1 U71 ( .A(n250), .Y(n194) );
  AND2X1 U72 ( .A(n218), .B(srstz), .Y(N298) );
  INVX1 U73 ( .A(n203), .Y(n211) );
  NAND21X1 U74 ( .B(n162), .A(n184), .Y(n174) );
  NAND32X1 U75 ( .B(n35), .C(n130), .A(n155), .Y(n99) );
  NAND21X1 U76 ( .B(n94), .A(n92), .Y(n51) );
  NAND21X1 U77 ( .B(n77), .A(n38), .Y(n42) );
  MUX2BXL U78 ( .D0(n82), .D1(n81), .S(n80), .Y(n83) );
  INVX1 U79 ( .A(n93), .Y(n80) );
  NAND21X1 U80 ( .B(n99), .A(n91), .Y(n81) );
  AO21X1 U81 ( .B(n51), .C(n42), .A(n57), .Y(n39) );
  AND3X1 U82 ( .A(n92), .B(n94), .C(n57), .Y(n59) );
  INVX1 U83 ( .A(n76), .Y(n92) );
  AND2X1 U84 ( .A(n205), .B(n206), .Y(ptx_crcshfo4) );
  NAND32X1 U85 ( .B(n57), .C(n76), .A(n79), .Y(n62) );
  NAND21X1 U86 ( .B(n203), .A(n161), .Y(n184) );
  INVX1 U87 ( .A(n31), .Y(n37) );
  AND2X1 U88 ( .A(n216), .B(srstz), .Y(N299) );
  INVX1 U89 ( .A(n65), .Y(n89) );
  INVX1 U90 ( .A(n103), .Y(n112) );
  INVX1 U91 ( .A(n172), .Y(n205) );
  INVX1 U92 ( .A(n216), .Y(n219) );
  NAND21X1 U93 ( .B(ptx_crcsidat[3]), .A(n32), .Y(n21) );
  NAND21X1 U94 ( .B(n187), .A(n199), .Y(n203) );
  NAND21X1 U95 ( .B(n187), .A(n5), .Y(n143) );
  NAND21X1 U96 ( .B(n2), .A(n221), .Y(ptx_fifopop) );
  AND4X1 U97 ( .A(r_txnumk[2]), .B(r_txnumk[3]), .C(r_txnumk[1]), .D(
        r_txnumk[0]), .Y(n26) );
  INVX3 U98 ( .A(n215), .Y(n77) );
  INVX1 U99 ( .A(i_rdat[5]), .Y(n127) );
  INVX1 U100 ( .A(i_rdat[3]), .Y(n152) );
  INVX1 U101 ( .A(i_rdat[2]), .Y(n153) );
  INVX1 U102 ( .A(i_one), .Y(n139) );
  INVX1 U103 ( .A(n207), .Y(n25) );
  INVX1 U104 ( .A(n214), .Y(n23) );
  INVX1 U105 ( .A(n175), .Y(n145) );
  INVX1 U106 ( .A(n125), .Y(n151) );
  NAND21XL U107 ( .B(i_rdat[6]), .A(n124), .Y(n125) );
  NAND21X1 U108 ( .B(n146), .A(prx_cccnt[0]), .Y(n187) );
  INVX1 U109 ( .A(ptx_txact), .Y(n146) );
  NAND32X1 U110 ( .B(n176), .C(n159), .A(n170), .Y(n155) );
  INVX1 U111 ( .A(n217), .Y(n210) );
  AO21X1 U112 ( .B(n242), .C(n193), .A(N252), .Y(n195) );
  AOI21BX1 U113 ( .C(n227), .B(n8), .A(n174), .Y(n179) );
  AOI21X1 U114 ( .B(n245), .C(n244), .A(ptx_txact), .Y(n8) );
  OAI211X1 U115 ( .C(n160), .D(n159), .A(n158), .B(n157), .Y(n218) );
  AOI221XL U116 ( .A(n205), .B(n171), .C(n210), .D(n173), .E(n142), .Y(n160)
         );
  OA22X1 U117 ( .A(n173), .B(n156), .C(n162), .D(n155), .Y(n157) );
  AOI32X1 U118 ( .A(i_txreq), .B(n244), .C(n146), .D(n145), .E(n144), .Y(n158)
         );
  INVX1 U119 ( .A(n202), .Y(n220) );
  NAND21X1 U120 ( .B(n190), .A(n193), .Y(n250) );
  AND4XL U121 ( .A(n215), .B(n214), .C(n213), .D(n212), .Y(ptx_crcstart) );
  AND2X1 U122 ( .A(srstz), .B(n202), .Y(N297) );
  AND3XL U123 ( .A(n210), .B(n215), .C(n206), .Y(ptx_crcshfi4) );
  NAND32X1 U124 ( .B(n169), .C(n174), .A(n168), .Y(n216) );
  INVX1 U125 ( .A(n173), .Y(n169) );
  AO21X1 U126 ( .B(n177), .C(n172), .A(n170), .Y(n168) );
  INVX1 U127 ( .A(n221), .Y(n162) );
  INVX1 U128 ( .A(n167), .Y(n177) );
  OAI31XL U129 ( .A(n166), .B(n165), .C(n175), .D(n164), .Y(n167) );
  INVX1 U130 ( .A(n163), .Y(n166) );
  INVX1 U131 ( .A(n164), .Y(n142) );
  NAND21X1 U132 ( .B(n98), .A(n38), .Y(n76) );
  MUX2X1 U133 ( .D0(n224), .D1(n120), .S(n119), .Y(n121) );
  XOR2X1 U134 ( .A(n192), .B(n118), .Y(n119) );
  MUX3X1 U135 ( .D0(n116), .D1(n115), .D2(n114), .S0(n113), .S1(n17), .Y(n120)
         );
  MUX4X1 U136 ( .D0(encout[0]), .D1(encout[1]), .D2(encout[2]), .D3(encout[3]), 
        .S0(n17), .S1(N45), .Y(n224) );
  NAND43X1 U137 ( .B(n161), .C(n110), .D(n86), .A(n85), .Y(encout[3]) );
  OAI32XL U138 ( .A(n77), .B(n79), .C(n76), .D(n75), .E(n155), .Y(n86) );
  AOI221XL U139 ( .A(i_rdat[3]), .B(n112), .C(n95), .D(n84), .E(n83), .Y(n85)
         );
  AND3X1 U140 ( .A(n74), .B(n73), .C(n72), .Y(n75) );
  AO21X1 U141 ( .B(n112), .C(n111), .A(n110), .Y(n114) );
  MUX2XL U142 ( .D0(i_rdat[7]), .D1(i_rdat[5]), .S(n113), .Y(n111) );
  NAND21X1 U143 ( .B(n165), .A(n163), .Y(n144) );
  INVX1 U144 ( .A(N45), .Y(n113) );
  OAI221X1 U145 ( .A(n76), .B(n100), .C(n103), .D(n150), .E(n39), .Y(n41) );
  NAND21X1 U146 ( .B(n235), .A(n43), .Y(n40) );
  NAND5XL U147 ( .A(n65), .B(n64), .C(n63), .D(n62), .E(n61), .Y(encout[2]) );
  AOI221XL U148 ( .A(n79), .B(n95), .C(i_rdat[2]), .D(n112), .E(n60), .Y(n61)
         );
  MUX2BXL U149 ( .D0(n59), .D1(n58), .S(n77), .Y(n60) );
  NAND21X1 U150 ( .B(n57), .A(n82), .Y(n58) );
  INVX1 U151 ( .A(n171), .Y(n165) );
  GEN2XL U152 ( .D(n94), .E(n98), .C(n48), .B(n95), .A(n47), .Y(n49) );
  OA21X1 U153 ( .B(n57), .C(n98), .A(n90), .Y(n48) );
  INVX1 U154 ( .A(n63), .Y(n47) );
  NAND43X1 U155 ( .B(n109), .C(n108), .D(n107), .A(n106), .Y(n115) );
  INVX1 U156 ( .A(n105), .Y(n106) );
  AND3X1 U157 ( .A(n92), .B(n91), .C(n90), .Y(n109) );
  AND3X1 U158 ( .A(n95), .B(n94), .C(n93), .Y(n108) );
  NAND21X1 U159 ( .B(n56), .A(n55), .Y(encout[1]) );
  AOI211X1 U160 ( .C(n54), .D(n91), .A(n53), .B(n110), .Y(n55) );
  OA21XL U161 ( .B(n215), .C(n90), .A(n82), .Y(n53) );
  AOI211X1 U162 ( .C(n231), .D(n223), .A(n97), .B(n96), .Y(n104) );
  AO21X1 U163 ( .B(n101), .C(n100), .A(n99), .Y(n102) );
  INVX1 U164 ( .A(n229), .Y(n96) );
  AO21XL U165 ( .B(i_rdat[6]), .C(n112), .A(n89), .Y(n116) );
  INVX1 U166 ( .A(n84), .Y(n94) );
  INVX1 U167 ( .A(n78), .Y(n57) );
  NAND31X1 U168 ( .C(n145), .A(n9), .B(n65), .Y(n110) );
  NAND21X1 U169 ( .B(n79), .A(n78), .Y(n93) );
  AO21X1 U170 ( .B(n242), .C(n190), .A(n117), .Y(n118) );
  NAND32XL U171 ( .B(n215), .C(n78), .A(n79), .Y(n100) );
  INVX1 U172 ( .A(n90), .Y(n79) );
  OA21X1 U173 ( .B(n223), .C(n228), .A(n235), .Y(n45) );
  INVX1 U174 ( .A(n98), .Y(n101) );
  INVX1 U175 ( .A(n50), .Y(n91) );
  NAND21XL U176 ( .B(n215), .A(n94), .Y(n50) );
  INVX1 U177 ( .A(n97), .Y(n74) );
  NAND32X1 U178 ( .B(n170), .C(n159), .A(n176), .Y(n172) );
  INVX1 U179 ( .A(n222), .Y(ptx_goidle) );
  INVX1 U180 ( .A(n140), .Y(n35) );
  INVX1 U181 ( .A(r_txauto[4]), .Y(n156) );
  INVX1 U182 ( .A(n64), .Y(n161) );
  AND4X1 U183 ( .A(n220), .B(n219), .C(n218), .D(n217), .Y(ptx_pspyld) );
  AOI32X1 U184 ( .A(n208), .B(n28), .C(n209), .D(r_txnumk[4]), .E(n27), .Y(n29) );
  NAND21X1 U185 ( .B(n26), .A(bytcnt[4]), .Y(n27) );
  OAI31XL U186 ( .A(n25), .B(n24), .C(n23), .D(n22), .Y(n28) );
  MUX2X1 U187 ( .D0(n154), .D1(n127), .S(hinib), .Y(n36) );
  INVX1 U188 ( .A(bytcnt[3]), .Y(n136) );
  INVX1 U189 ( .A(bytcnt[2]), .Y(n135) );
  INVX1 U190 ( .A(bytcnt[4]), .Y(n134) );
  AOI22BX1 U191 ( .B(bytcnt[0]), .A(r_txnumk[0]), .D(bytcnt[1]), .C(
        r_txnumk[1]), .Y(n24) );
  NAND21X1 U192 ( .B(r_txnumk[4]), .A(bytcnt[4]), .Y(n208) );
  NAND21XL U193 ( .B(r_txnumk[3]), .A(bytcnt[3]), .Y(n209) );
  NAND21X1 U194 ( .B(n139), .A(r_txendk), .Y(n148) );
  INVX1 U195 ( .A(n129), .Y(n199) );
  XOR2X1 U196 ( .A(n130), .B(bitcnt[2]), .Y(n132) );
  NAND32X1 U197 ( .B(ptx_fsm[0]), .C(n159), .A(n170), .Y(n217) );
  INVX1 U198 ( .A(ptx_fsm[1]), .Y(n159) );
  NAND32X1 U199 ( .B(ptx_fsm[1]), .C(n176), .A(n170), .Y(n175) );
  INVX1 U200 ( .A(ptx_fsm[2]), .Y(n170) );
  INVX1 U201 ( .A(ptx_fsm[0]), .Y(n176) );
  OR2X1 U202 ( .A(ptx_fsm[2]), .B(n198), .Y(ptx_txact) );
  NAND21X1 U203 ( .B(ptx_fsm[1]), .A(n176), .Y(n198) );
  INVX1 U204 ( .A(bitcnt[0]), .Y(n190) );
  AND3X1 U205 ( .A(n12), .B(n13), .C(n181), .Y(n11) );
  XNOR2XL U206 ( .A(n218), .B(ptx_fsm[1]), .Y(n12) );
  AOI21X1 U207 ( .B(n216), .C(n170), .A(i_txreq), .Y(n13) );
  OAI211X1 U208 ( .C(r_txauto[5]), .D(n180), .A(n179), .B(n178), .Y(n202) );
  OA22X1 U209 ( .A(r_txauto[4]), .B(n173), .C(n172), .D(n171), .Y(n180) );
  OA22X1 U210 ( .A(n177), .B(n176), .C(n245), .D(n175), .Y(n178) );
  XOR2X1 U211 ( .A(ptx_fsm[0]), .B(n220), .Y(n181) );
  MUX2IX1 U212 ( .D0(n14), .D1(n15), .S(bitcnt[3]), .Y(N255) );
  NAND3X1 U213 ( .A(bitcnt[2]), .B(n194), .C(bitcnt[1]), .Y(n14) );
  AOI21X1 U214 ( .B(n193), .C(n192), .A(n195), .Y(n15) );
  NAND5XL U215 ( .A(bytcnt[1]), .B(bytcnt[0]), .C(bytcnt[2]), .D(bytcnt[3]), 
        .E(bytcnt[4]), .Y(n182) );
  AOI31XL U216 ( .A(n155), .B(n175), .C(n172), .D(n143), .Y(n183) );
  INVX1 U217 ( .A(n189), .Y(N252) );
  NAND21X1 U218 ( .B(bitcnt[0]), .A(n193), .Y(n189) );
  MUX2X1 U219 ( .D0(n196), .D1(n195), .S(bitcnt[2]), .Y(N254) );
  AND2X1 U220 ( .A(n194), .B(bitcnt[1]), .Y(n196) );
  MUX2IX1 U221 ( .D0(n226), .D1(n225), .S(n16), .Y(n238) );
  NAND3X1 U222 ( .A(srstz), .B(n227), .C(n123), .Y(n16) );
  AOI211XL U223 ( .C(n199), .D(n198), .A(i_txreq), .B(n5), .Y(n200) );
  OAI31XL U224 ( .A(n155), .B(bytcnt[1]), .C(n147), .D(n141), .Y(n164) );
  AND4X1 U225 ( .A(n217), .B(n222), .C(n172), .D(n175), .Y(n141) );
  NAND21XL U226 ( .B(n143), .A(r_txshrt), .Y(n163) );
  NAND21X1 U227 ( .B(n138), .A(n137), .Y(n171) );
  INVXL U228 ( .A(n147), .Y(n137) );
  MUX2X1 U229 ( .D0(n187), .D1(n122), .S(prx_cccnt[1]), .Y(n123) );
  NAND21X1 U230 ( .B(n146), .A(n121), .Y(n122) );
  NAND21X1 U231 ( .B(n190), .A(n87), .Y(n88) );
  INVXL U232 ( .A(n130), .Y(n87) );
  GEN2XL U233 ( .D(n1), .E(n231), .C(n34), .B(n33), .A(n89), .Y(n105) );
  INVX1 U234 ( .A(n155), .Y(n33) );
  INVX1 U235 ( .A(n73), .Y(n34) );
  MUX2X1 U236 ( .D0(ptx_crcsidat[0]), .D1(pcc_crc30[0]), .S(n205), .Y(n78) );
  MUX2XL U237 ( .D0(ptx_crcsidat[3]), .D1(pcc_crc30[3]), .S(n205), .Y(n98) );
  MUX2XL U238 ( .D0(ptx_crcsidat[2]), .D1(pcc_crc30[2]), .S(n205), .Y(n84) );
  NAND21XL U239 ( .B(n130), .A(n1), .Y(n117) );
  XNOR2XL U240 ( .A(n117), .B(bitcnt[0]), .Y(n17) );
  MUX2BXL U241 ( .D0(n36), .D1(pcc_crc30[1]), .S(n205), .Y(n90) );
  NAND21X1 U242 ( .B(n155), .A(n46), .Y(n63) );
  MUX2X1 U243 ( .D0(n223), .D1(n43), .S(r_txauto[0]), .Y(n44) );
  OAI221X1 U244 ( .A(n232), .B(n71), .C(n70), .D(n240), .E(n69), .Y(n97) );
  INVX1 U245 ( .A(n234), .Y(n70) );
  NAND21X1 U246 ( .B(n230), .A(n66), .Y(n67) );
  NAND21X1 U247 ( .B(n233), .A(n223), .Y(n68) );
  INVX1 U248 ( .A(n235), .Y(n66) );
  INVX1 U249 ( .A(n233), .Y(n20) );
  NAND43X1 U250 ( .B(ptx_cc), .C(n187), .D(n140), .A(ptx_fsm[0]), .Y(n222) );
  NAND21X1 U251 ( .B(ptx_fsm[1]), .A(ptx_fsm[2]), .Y(n140) );
  NAND21X1 U252 ( .B(ptx_fsm[0]), .A(n35), .Y(n64) );
  INVX1 U253 ( .A(bitcnt[2]), .Y(n192) );
  XOR2X1 U254 ( .A(add_104_carry[4]), .B(bytcnt[4]), .Y(N267) );
  NOR2X1 U255 ( .A(n18), .B(n226), .Y(n225) );
  INVX1 U256 ( .A(ptx_cc), .Y(n226) );
  MUX2IX1 U257 ( .D0(n234), .D1(n239), .S(n230), .Y(n236) );
  INVX1 U258 ( .A(n240), .Y(n230) );
  NAND2X1 U259 ( .A(n235), .B(n233), .Y(n239) );
  INVX1 U260 ( .A(n228), .Y(n231) );
  AOI21BBXL U261 ( .B(n229), .C(n240), .A(n234), .Y(n241) );
  NOR21XL U262 ( .B(N267), .A(n243), .Y(N273) );
  NOR21XL U263 ( .B(N266), .A(n243), .Y(N272) );
  NOR21XL U264 ( .B(N265), .A(n243), .Y(N271) );
  NOR21XL U265 ( .B(N264), .A(n243), .Y(N270) );
  NOR21XL U266 ( .B(n223), .A(n243), .Y(N269) );
  NAND2X1 U267 ( .A(n11), .B(n243), .Y(N268) );
  NOR43XL U268 ( .B(n235), .C(n246), .D(n228), .A(n234), .Y(n245) );
  NOR3XL U269 ( .A(n247), .B(r_txauto[0]), .C(n248), .Y(n234) );
  NAND3X1 U270 ( .A(r_txauto[0]), .B(n248), .C(r_txauto[2]), .Y(n228) );
  AND3X1 U271 ( .A(n232), .B(n229), .C(n233), .Y(n246) );
  NAND3X1 U272 ( .A(n249), .B(n248), .C(r_txauto[2]), .Y(n233) );
  INVX1 U273 ( .A(r_txauto[0]), .Y(n249) );
  NAND3X1 U274 ( .A(n248), .B(n247), .C(r_txauto[0]), .Y(n229) );
  INVX1 U275 ( .A(r_txauto[1]), .Y(n248) );
  NAND2X1 U276 ( .A(r_txauto[1]), .B(n247), .Y(n232) );
  INVX1 U277 ( .A(r_txauto[2]), .Y(n247) );
  NAND3X1 U278 ( .A(r_txauto[2]), .B(r_txauto[0]), .C(r_txauto[1]), .Y(n235)
         );
  INVX1 U279 ( .A(r_txauto[3]), .Y(n244) );
  INVX1 U280 ( .A(i_txreq), .Y(n227) );
  MUX2BXL U281 ( .D0(N252), .D1(n250), .S(n242), .Y(N253) );
  INVX1 U282 ( .A(bitcnt[1]), .Y(n242) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phytx_a0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phytx_a0_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module phyidd_a0 ( i_trans, i_goidle, o_ccidle, o_goidle, o_gobusy, clk, srstz
 );
  input i_trans, i_goidle, clk, srstz;
  output o_ccidle, o_goidle, o_gobusy;
  wire   N11, N12, N13, N14, N15, N16, N17, N18, N46, N47, N48, N49, N50, N51,
         N52, N53, N55, N56, N57, N58, N59, N60, N61, N62, N73, N74, N75, N76,
         N77, N78, N79, N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N90,
         N91, net10611, net10617, net10622, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27;
  wire   [7:0] ttranwin;
  wire   [1:0] ntrancnt;
  wire   [7:0] trans0;
  wire   [7:0] ttranwin_minus;
  wire   [7:0] trans1;

  SNPS_CLOCK_GATE_HIGH_phyidd_a0_0 clk_gate_trans1_reg ( .CLK(clk), .EN(N90), 
        .ENCLK(net10611), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_phyidd_a0_2 clk_gate_trans0_reg ( .CLK(clk), .EN(N91), 
        .ENCLK(net10617), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_phyidd_a0_1 clk_gate_ttranwin_reg ( .CLK(clk), .EN(N81), 
        .ENCLK(net10622), .TE(1'b0) );
  phyidd_a0_DW01_sub_0 sub_47 ( .A(trans1), .B(trans0), .CI(1'b0), .DIFF({N53, 
        N52, N51, N50, N49, N48, N47, N46}), .CO() );
  phyidd_a0_DW01_sub_1 sub_24 ( .A({n27, n26, n25, n24, n23, n22, n21, n20}), 
        .B(trans0), .CI(1'b0), .DIFF(ttranwin_minus), .CO() );
  phyidd_a0_DW01_inc_0 add_23 ( .A(ttranwin), .SUM({N18, N17, N16, N15, N14, 
        N13, N12, N11}) );
  DFFQX1 trans1_reg_6_ ( .D(N79), .C(net10611), .Q(trans1[6]) );
  DFFQX1 trans1_reg_7_ ( .D(N80), .C(net10611), .Q(trans1[7]) );
  DFFQX1 trans0_reg_7_ ( .D(N62), .C(net10617), .Q(trans0[7]) );
  DFFQX1 trans1_reg_4_ ( .D(N77), .C(net10611), .Q(trans1[4]) );
  DFFQX1 trans1_reg_5_ ( .D(N78), .C(net10611), .Q(trans1[5]) );
  DFFQX1 trans0_reg_5_ ( .D(N60), .C(net10617), .Q(trans0[5]) );
  DFFQX1 trans0_reg_6_ ( .D(N61), .C(net10617), .Q(trans0[6]) );
  DFFQX1 trans1_reg_3_ ( .D(N76), .C(net10611), .Q(trans1[3]) );
  DFFQX1 ntrancnt_reg_1_ ( .D(n56), .C(clk), .Q(ntrancnt[1]) );
  DFFQX1 ntrancnt_reg_0_ ( .D(n57), .C(clk), .Q(ntrancnt[0]) );
  DFFQX1 trans0_reg_4_ ( .D(N59), .C(net10617), .Q(trans0[4]) );
  DFFQX1 trans1_reg_1_ ( .D(N74), .C(net10611), .Q(trans1[1]) );
  DFFQX1 trans1_reg_2_ ( .D(N75), .C(net10611), .Q(trans1[2]) );
  DFFQX1 trans0_reg_2_ ( .D(N57), .C(net10617), .Q(trans0[2]) );
  DFFQX1 trans0_reg_3_ ( .D(N58), .C(net10617), .Q(trans0[3]) );
  DFFQX1 trans1_reg_0_ ( .D(N73), .C(net10611), .Q(trans1[0]) );
  DFFQX1 trans0_reg_0_ ( .D(N55), .C(net10617), .Q(trans0[0]) );
  DFFQX1 trans0_reg_1_ ( .D(N56), .C(net10617), .Q(trans0[1]) );
  DFFQX1 ttranwin_reg_7_ ( .D(N89), .C(net10622), .Q(ttranwin[7]) );
  DFFQX1 ttranwin_reg_5_ ( .D(N87), .C(net10622), .Q(ttranwin[5]) );
  DFFQX1 ttranwin_reg_1_ ( .D(N83), .C(net10622), .Q(ttranwin[1]) );
  DFFQX1 ttranwin_reg_6_ ( .D(N88), .C(net10622), .Q(ttranwin[6]) );
  DFFQX1 ttranwin_reg_0_ ( .D(N82), .C(net10622), .Q(ttranwin[0]) );
  DFFQX1 ttranwin_reg_4_ ( .D(N86), .C(net10622), .Q(ttranwin[4]) );
  DFFQX1 ttranwin_reg_2_ ( .D(N84), .C(net10622), .Q(ttranwin[2]) );
  DFFQX1 ttranwin_reg_3_ ( .D(N85), .C(net10622), .Q(ttranwin[3]) );
  DFFQX1 ccidle_reg ( .D(n55), .C(clk), .Q(o_ccidle) );
  NAND2X1 U3 ( .A(ntrancnt[0]), .B(n18), .Y(n3) );
  NAND2X1 U4 ( .A(ntrancnt[1]), .B(n16), .Y(n4) );
  INVX1 U5 ( .A(n37), .Y(o_goidle) );
  OAI22X1 U6 ( .A(n30), .B(n47), .C(n46), .D(n6), .Y(N88) );
  OAI22X1 U7 ( .A(n31), .B(n47), .C(n46), .D(n7), .Y(N87) );
  OAI22X1 U8 ( .A(n32), .B(n47), .C(n46), .D(n8), .Y(N86) );
  NAND2X1 U11 ( .A(n50), .B(n17), .Y(n46) );
  OAI22X1 U12 ( .A(n33), .B(n47), .C(n46), .D(n9), .Y(N85) );
  OAI22X1 U13 ( .A(n34), .B(n47), .C(n46), .D(n10), .Y(N84) );
  OAI22X1 U14 ( .A(n35), .B(n47), .C(n46), .D(n11), .Y(N83) );
  INVX1 U15 ( .A(n50), .Y(n13) );
  NAND2X1 U16 ( .A(N12), .B(n45), .Y(n35) );
  INVX1 U17 ( .A(n36), .Y(n20) );
  OAI22X1 U18 ( .A(n29), .B(n41), .C(n43), .D(n5), .Y(N80) );
  OAI22X1 U19 ( .A(n29), .B(n47), .C(n46), .D(n5), .Y(N89) );
  AOI21X1 U20 ( .B(n15), .C(n19), .A(i_goidle), .Y(n37) );
  INVX1 U21 ( .A(ttranwin_minus[6]), .Y(n6) );
  NAND2X1 U22 ( .A(N13), .B(n45), .Y(n34) );
  OAI22X1 U23 ( .A(n30), .B(n4), .C(n43), .D(n6), .Y(N79) );
  NOR3XL U24 ( .A(n14), .B(n41), .C(n19), .Y(o_gobusy) );
  INVX1 U25 ( .A(ttranwin_minus[5]), .Y(n7) );
  INVX1 U26 ( .A(ttranwin_minus[4]), .Y(n8) );
  NAND2X1 U27 ( .A(N14), .B(n45), .Y(n33) );
  NAND2X1 U28 ( .A(N15), .B(n45), .Y(n32) );
  OAI222XL U29 ( .A(n38), .B(n18), .C(n39), .D(n3), .E(n41), .F(n39), .Y(n56)
         );
  INVX1 U30 ( .A(i_trans), .Y(n14) );
  EORX1 U31 ( .A(n39), .B(n42), .C(n39), .D(n43), .Y(n38) );
  OAI22X1 U32 ( .A(n31), .B(n41), .C(n43), .D(n7), .Y(N78) );
  OAI22X1 U33 ( .A(n32), .B(n4), .C(n43), .D(n8), .Y(N77) );
  NAND2X1 U34 ( .A(n42), .B(i_trans), .Y(n39) );
  NOR3XL U35 ( .A(o_gobusy), .B(o_goidle), .C(n44), .Y(n42) );
  OAI21X1 U36 ( .B(n45), .C(i_trans), .A(srstz), .Y(n44) );
  NAND31X1 U37 ( .C(N91), .A(n48), .B(n51), .Y(N81) );
  AOI21BBXL U38 ( .B(n13), .C(n4), .A(n52), .Y(n51) );
  NAND32X1 U39 ( .B(n52), .C(n15), .A(n14), .Y(n48) );
  AND2X1 U40 ( .A(n48), .B(n49), .Y(n47) );
  OAI21BBX1 U41 ( .A(n4), .B(n40), .C(n50), .Y(n49) );
  INVX1 U42 ( .A(ttranwin_minus[3]), .Y(n9) );
  NOR2X1 U43 ( .A(n52), .B(n14), .Y(n50) );
  NOR2X1 U44 ( .A(n15), .B(N17), .Y(n30) );
  NAND2X1 U45 ( .A(N16), .B(n45), .Y(n31) );
  OAI21X1 U46 ( .B(n40), .C(n13), .A(n46), .Y(N91) );
  OAI22X1 U47 ( .A(n36), .B(n47), .C(n46), .D(n12), .Y(N82) );
  OAI22X1 U48 ( .A(n33), .B(n41), .C(n43), .D(n9), .Y(N76) );
  ENOX1 U49 ( .A(n30), .B(n3), .C(N52), .D(n17), .Y(N61) );
  ENOX1 U50 ( .A(n31), .B(n40), .C(N51), .D(n17), .Y(N60) );
  INVX1 U51 ( .A(n45), .Y(n15) );
  INVX1 U52 ( .A(ttranwin_minus[2]), .Y(n10) );
  INVX1 U53 ( .A(ttranwin_minus[1]), .Y(n11) );
  OAI22X1 U54 ( .A(n34), .B(n4), .C(n43), .D(n10), .Y(N75) );
  OAI22X1 U55 ( .A(n35), .B(n41), .C(n43), .D(n11), .Y(N74) );
  OAI21X1 U56 ( .B(n41), .C(n13), .A(n46), .Y(N90) );
  ENOX1 U57 ( .A(n32), .B(n3), .C(N50), .D(n17), .Y(N59) );
  OAI211X1 U58 ( .C(o_gobusy), .D(n19), .A(n37), .B(srstz), .Y(n55) );
  INVX1 U59 ( .A(ttranwin_minus[0]), .Y(n12) );
  OAI22X1 U60 ( .A(n36), .B(n4), .C(n43), .D(n12), .Y(N73) );
  ENOX1 U61 ( .A(n33), .B(n40), .C(N49), .D(n17), .Y(N58) );
  ENOX1 U62 ( .A(n34), .B(n3), .C(N48), .D(n17), .Y(N57) );
  INVX1 U63 ( .A(n43), .Y(n17) );
  ENOX1 U64 ( .A(n35), .B(n40), .C(N47), .D(n17), .Y(N56) );
  INVX1 U65 ( .A(n34), .Y(n22) );
  INVX1 U66 ( .A(n33), .Y(n23) );
  INVX1 U67 ( .A(n32), .Y(n24) );
  INVX1 U68 ( .A(n31), .Y(n25) );
  INVX1 U69 ( .A(n30), .Y(n26) );
  NAND4X1 U70 ( .A(ttranwin[7]), .B(ttranwin[6]), .C(n53), .D(n54), .Y(n45) );
  NOR2X1 U71 ( .A(ttranwin[1]), .B(ttranwin[0]), .Y(n53) );
  NOR4XL U72 ( .A(ttranwin[5]), .B(ttranwin[4]), .C(ttranwin[3]), .D(
        ttranwin[2]), .Y(n54) );
  INVX1 U73 ( .A(n35), .Y(n21) );
  INVX1 U74 ( .A(ttranwin_minus[7]), .Y(n5) );
  INVX1 U75 ( .A(n29), .Y(n27) );
  NAND2X1 U76 ( .A(N11), .B(n45), .Y(n36) );
  ENOX1 U77 ( .A(n29), .B(n3), .C(N53), .D(n17), .Y(N62) );
  OAI31XL U78 ( .A(n19), .B(ntrancnt[0]), .C(n14), .D(srstz), .Y(n52) );
  NOR2X1 U79 ( .A(n15), .B(N18), .Y(n29) );
  OAI22X1 U80 ( .A(n38), .B(n16), .C(ntrancnt[0]), .D(n39), .Y(n57) );
  INVX1 U81 ( .A(o_ccidle), .Y(n19) );
  NAND2X1 U82 ( .A(ntrancnt[1]), .B(n16), .Y(n41) );
  INVX1 U83 ( .A(ntrancnt[0]), .Y(n16) );
  NAND2X1 U84 ( .A(ntrancnt[0]), .B(ntrancnt[1]), .Y(n43) );
  NAND2X1 U85 ( .A(ntrancnt[0]), .B(n18), .Y(n40) );
  INVX1 U86 ( .A(ntrancnt[1]), .Y(n18) );
  ENOX1 U87 ( .A(n36), .B(n40), .C(N46), .D(n17), .Y(N55) );
endmodule


module phyidd_a0_DW01_inc_0 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  XOR2X1 U1 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module phyidd_a0_DW01_sub_1 ( A, B, CI, DIFF, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9;
  wire   [7:1] carry;

  FAD1X1 U2_6 ( .A(A[6]), .B(n9), .CI(carry[6]), .CO(carry[7]), .SO(DIFF[6])
         );
  FAD1X1 U2_5 ( .A(A[5]), .B(n8), .CI(carry[5]), .CO(carry[6]), .SO(DIFF[5])
         );
  FAD1X1 U2_4 ( .A(A[4]), .B(n7), .CI(carry[4]), .CO(carry[5]), .SO(DIFF[4])
         );
  FAD1X1 U2_3 ( .A(A[3]), .B(n6), .CI(carry[3]), .CO(carry[4]), .SO(DIFF[3])
         );
  FAD1X1 U2_2 ( .A(A[2]), .B(n5), .CI(carry[2]), .CO(carry[3]), .SO(DIFF[2])
         );
  FAD1X1 U2_1 ( .A(A[1]), .B(n4), .CI(carry[1]), .CO(carry[2]), .SO(DIFF[1])
         );
  XOR3X1 U2_7 ( .A(A[7]), .B(n3), .C(carry[7]), .Y(DIFF[7]) );
  INVX1 U1 ( .A(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(DIFF[0]) );
  INVX1 U3 ( .A(B[2]), .Y(n5) );
  INVX1 U4 ( .A(B[3]), .Y(n6) );
  INVX1 U5 ( .A(B[4]), .Y(n7) );
  INVX1 U6 ( .A(B[5]), .Y(n8) );
  INVX1 U7 ( .A(B[6]), .Y(n9) );
  INVX1 U8 ( .A(B[1]), .Y(n4) );
  NAND21X1 U9 ( .B(n2), .A(n1), .Y(carry[1]) );
  INVX1 U10 ( .A(B[7]), .Y(n3) );
  INVX1 U11 ( .A(B[0]), .Y(n2) );
endmodule


module phyidd_a0_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9;
  wire   [7:1] carry;

  FAD1X1 U2_6 ( .A(A[6]), .B(n9), .CI(carry[6]), .CO(carry[7]), .SO(DIFF[6])
         );
  FAD1X1 U2_5 ( .A(A[5]), .B(n8), .CI(carry[5]), .CO(carry[6]), .SO(DIFF[5])
         );
  FAD1X1 U2_4 ( .A(A[4]), .B(n7), .CI(carry[4]), .CO(carry[5]), .SO(DIFF[4])
         );
  FAD1X1 U2_3 ( .A(A[3]), .B(n6), .CI(carry[3]), .CO(carry[4]), .SO(DIFF[3])
         );
  FAD1X1 U2_2 ( .A(A[2]), .B(n5), .CI(carry[2]), .CO(carry[3]), .SO(DIFF[2])
         );
  FAD1X1 U2_1 ( .A(A[1]), .B(n4), .CI(carry[1]), .CO(carry[2]), .SO(DIFF[1])
         );
  XOR3X1 U2_7 ( .A(A[7]), .B(n3), .C(carry[7]), .Y(DIFF[7]) );
  INVX1 U1 ( .A(B[2]), .Y(n5) );
  INVX1 U2 ( .A(B[3]), .Y(n6) );
  INVX1 U3 ( .A(B[4]), .Y(n7) );
  INVX1 U4 ( .A(B[5]), .Y(n8) );
  INVX1 U5 ( .A(B[6]), .Y(n9) );
  INVX1 U6 ( .A(B[1]), .Y(n4) );
  NAND21X1 U7 ( .B(n2), .A(n1), .Y(carry[1]) );
  INVX1 U8 ( .A(A[0]), .Y(n1) );
  INVX1 U9 ( .A(B[0]), .Y(n2) );
  INVX1 U10 ( .A(B[7]), .Y(n3) );
  XOR2X1 U11 ( .A(B[0]), .B(A[0]), .Y(DIFF[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyidd_a0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyidd_a0_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyidd_a0_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module phyrx_a0 ( i_cc, ptx_txact, r_adprx_en, r_adp2nd, r_exist1st, r_ordrs4, 
        r_rxdb_opt, r_ords_ena, r_pshords, r_rgdcrc, prx_cccnt, prx_rst, 
        prx_setsta, prx_idle, prx_d_cc, prx_bmc, prx_trans, prx_fiforst, 
        prx_fifopsh, prx_fifowdat, pff_txreq, pid_gobusy, pid_goidle, 
        pid_ccidle, pcc_rxgood, prx_crcstart, prx_crcshfi4, prx_crcsidat, 
        prx_rxcode, prx_adpn, prx_rcvdords, prx_eoprcvd, prx_fsm, clk, srstz
 );
  input [1:0] r_rxdb_opt;
  input [6:0] r_ords_ena;
  output [1:0] prx_cccnt;
  output [1:0] prx_rst;
  output [6:0] prx_setsta;
  output [7:0] prx_fifowdat;
  output [3:0] prx_crcsidat;
  output [4:0] prx_rxcode;
  output [5:0] prx_adpn;
  output [2:0] prx_rcvdords;
  output [3:0] prx_fsm;
  input i_cc, ptx_txact, r_adprx_en, r_adp2nd, r_exist1st, r_ordrs4, r_pshords,
         r_rgdcrc, pff_txreq, pid_gobusy, pid_goidle, pid_ccidle, pcc_rxgood,
         clk, srstz;
  output prx_idle, prx_d_cc, prx_bmc, prx_trans, prx_fiforst, prx_fifopsh,
         prx_crcstart, prx_crcshfi4, prx_eoprcvd;
  wire   N31, N32, N33, n267, n268, n269, db_gohi, db_golo, k0_det, cctrans,
         shrtrans, N58, N59, N60, N61, N62, N70, N71, N72, N73, N74, N75, N76,
         N96, N153, N154, N155, N156, N157, ps_ords_ena, cs_ords_ena, N236,
         N238, N239, N246, N247, N248, N249, N250, N251, N275, N276, N277,
         N278, N279, net10639, net10645, net10650, net10655, net10660,
         net10665, net10670, n21, n214, n1, n2, n3, n6, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n25, n28, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n263, n264, n265, n266;
  wire   [5:0] cccnt;
  wire   [2:0] ps_dat5b;
  wire   [2:0] bcnt;
  wire   [7:3] ordsbuf;
  wire   [5:2] add_83_carry;

  phyrx_db u0_phyrx_db ( .clk(clk), .srstz(srstz), .x_cc(i_cc), .ptx_txact(n8), 
        .r_rxdb_opt(r_rxdb_opt), .gohi(db_gohi), .golo(db_golo), .gotrans(
        prx_trans) );
  phyrx_adp u0_phyrx_adp ( .clk(clk), .srstz(srstz), .gohi(db_gohi), .golo(
        db_golo), .gobusy(pid_gobusy), .goidle(pid_goidle), .i_ccidle(
        pid_ccidle), .k0_det(k0_det), .r_adprx_en(r_adprx_en), .r_adp2nd(
        r_adp2nd), .adp_val(prx_adpn), .d_cc(prx_d_cc), .cctrans(cctrans) );
  SNPS_CLOCK_GATE_HIGH_phyrx_a0_0 clk_gate_cccnt_reg ( .CLK(clk), .EN(N70), 
        .ENCLK(net10639), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_phyrx_a0_6 clk_gate_cs_dat5b_reg ( .CLK(clk), .EN(N153), 
        .ENCLK(net10645), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_phyrx_a0_5 clk_gate_bcnt_reg ( .CLK(clk), .EN(N236), 
        .ENCLK(net10650), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_phyrx_a0_4 clk_gate_cs_dat4b_reg ( .CLK(clk), .EN(n21), 
        .ENCLK(net10655), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_phyrx_a0_3 clk_gate_ordsbuf_reg ( .CLK(clk), .EN(N251), 
        .ENCLK(net10660), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_phyrx_a0_2 clk_gate_ordsbuf_reg_0 ( .CLK(clk), .EN(N250), .ENCLK(net10665), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_phyrx_a0_1 clk_gate_cs_bmni_reg ( .CLK(clk), .EN(N275), 
        .ENCLK(net10670), .TE(1'b0) );
  HAD1X1 add_83_U1_1_1 ( .A(cccnt[1]), .B(cccnt[0]), .CO(add_83_carry[2]), 
        .SO(N58) );
  HAD1X1 add_83_U1_1_2 ( .A(cccnt[2]), .B(add_83_carry[2]), .CO(
        add_83_carry[3]), .SO(N59) );
  HAD1X1 add_83_U1_1_3 ( .A(cccnt[3]), .B(add_83_carry[3]), .CO(
        add_83_carry[4]), .SO(N60) );
  HAD1X1 add_83_U1_1_4 ( .A(cccnt[4]), .B(add_83_carry[4]), .CO(
        add_83_carry[5]), .SO(N61) );
  DFFQX1 cs_dat4b_reg_1_ ( .D(prx_crcsidat[1]), .C(net10655), .Q(
        prx_fifowdat[1]) );
  DFFQX1 ordsbuf_reg_3_ ( .D(N249), .C(net10665), .Q(ordsbuf[3]) );
  DFFQX1 ordsbuf_reg_4_ ( .D(prx_fifowdat[4]), .C(net10660), .Q(ordsbuf[4]) );
  DFFQX1 ordsbuf_reg_7_ ( .D(prx_fifowdat[7]), .C(net10660), .Q(ordsbuf[7]) );
  DFFQX1 ordsbuf_reg_6_ ( .D(prx_fifowdat[6]), .C(net10660), .Q(ordsbuf[6]) );
  DFFQX1 ordsbuf_reg_5_ ( .D(prx_fifowdat[5]), .C(net10660), .Q(ordsbuf[5]) );
  DFFQX1 cs_dat4b_reg_2_ ( .D(prx_fifowdat[6]), .C(net10655), .Q(n269) );
  DFFQX1 cs_dat4b_reg_0_ ( .D(prx_fifowdat[4]), .C(net10655), .Q(
        prx_fifowdat[0]) );
  DFFQX1 cs_dat4b_reg_3_ ( .D(prx_crcsidat[3]), .C(net10655), .Q(prx_rxcode[3]) );
  DFFQX1 cs_dat4b_reg_4_ ( .D(N96), .C(net10655), .Q(prx_rxcode[4]) );
  DFFQX1 bcnt_reg_1_ ( .D(N238), .C(net10650), .Q(bcnt[1]) );
  DFFQX1 bcnt_reg_2_ ( .D(N239), .C(net10650), .Q(bcnt[2]) );
  DFFQX1 bcnt_reg_0_ ( .D(n20), .C(net10650), .Q(bcnt[0]) );
  DFFQX1 cs_bmni_reg_1_ ( .D(N277), .C(net10670), .Q(prx_fsm[1]) );
  DFFQX1 cs_bmni_reg_2_ ( .D(N278), .C(net10670), .Q(prx_fsm[2]) );
  DFFQX1 cs_bmni_reg_0_ ( .D(N276), .C(net10670), .Q(prx_fsm[0]) );
  DFFQX1 cs_bmni_reg_3_ ( .D(N279), .C(net10670), .Q(prx_fsm[3]) );
  DFFQX1 cs_dat5b_reg_0_ ( .D(N154), .C(net10645), .Q(ps_dat5b[0]) );
  DFFQX1 cs_dat5b_reg_1_ ( .D(N155), .C(net10645), .Q(ps_dat5b[1]) );
  DFFQX1 cs_dat5b_reg_2_ ( .D(N156), .C(net10645), .Q(ps_dat5b[2]) );
  DFFQX1 cs_dat5b_reg_3_ ( .D(N157), .C(net10645), .Q(prx_bmc) );
  DFFQX1 cccnt_reg_4_ ( .D(N75), .C(net10639), .Q(cccnt[4]) );
  DFFQX1 shrtrans_reg ( .D(n214), .C(clk), .Q(shrtrans) );
  DFFQX1 cccnt_reg_5_ ( .D(N76), .C(net10639), .Q(cccnt[5]) );
  DFFQX1 cccnt_reg_1_ ( .D(N72), .C(net10639), .Q(cccnt[1]) );
  DFFQX1 cccnt_reg_3_ ( .D(N74), .C(net10639), .Q(cccnt[3]) );
  DFFQX1 cccnt_reg_2_ ( .D(N73), .C(net10639), .Q(cccnt[2]) );
  DFFQX1 cccnt_reg_0_ ( .D(N71), .C(net10639), .Q(cccnt[0]) );
  DFFQX1 ordsbuf_reg_2_ ( .D(N248), .C(net10665), .Q(prx_rcvdords[2]) );
  DFFQX1 ordsbuf_reg_1_ ( .D(N247), .C(net10665), .Q(prx_rcvdords[1]) );
  DFFQX1 ordsbuf_reg_0_ ( .D(N246), .C(net10665), .Q(prx_rcvdords[0]) );
  XOR2X1 U3 ( .A(n174), .B(ps_dat5b[2]), .Y(n49) );
  INVX3 U4 ( .A(n174), .Y(n148) );
  NAND31X4 U5 ( .C(n87), .A(cctrans), .B(n85), .Y(n174) );
  NAND21X1 U6 ( .B(n48), .A(prx_bmc), .Y(n41) );
  NAND2X1 U7 ( .A(n267), .B(prx_fifowdat[5]), .Y(n62) );
  INVX1 U8 ( .A(N96), .Y(n114) );
  NAND21X1 U9 ( .B(n58), .A(n53), .Y(n54) );
  AO21X1 U10 ( .B(n45), .C(n56), .A(n44), .Y(n46) );
  NAND21X1 U11 ( .B(n119), .A(n133), .Y(n120) );
  INVX1 U12 ( .A(n119), .Y(n21) );
  XNOR2XL U13 ( .A(prx_fsm[1]), .B(prx_fsm[0]), .Y(n1) );
  AOI21X1 U14 ( .B(n66), .C(n44), .A(n58), .Y(n2) );
  INVXL U15 ( .A(n269), .Y(n3) );
  INVXL U16 ( .A(n3), .Y(prx_fifowdat[2]) );
  INVX1 U17 ( .A(n115), .Y(prx_fifowdat[6]) );
  NAND21X1 U18 ( .B(n55), .A(n54), .Y(n267) );
  INVX1 U19 ( .A(n164), .Y(n6) );
  INVX1 U20 ( .A(n113), .Y(prx_fifowdat[4]) );
  NAND21X1 U21 ( .B(n47), .A(n46), .Y(n268) );
  BUFX3 U22 ( .A(ptx_txact), .Y(n8) );
  NAND32X1 U23 ( .B(n61), .C(n60), .A(n59), .Y(prx_fifowdat[5]) );
  BUFX3 U24 ( .A(prx_fifowdat[2]), .Y(prx_rxcode[2]) );
  BUFX3 U25 ( .A(prx_fifowdat[0]), .Y(prx_rxcode[0]) );
  BUFX3 U26 ( .A(prx_fifowdat[1]), .Y(prx_rxcode[1]) );
  NOR2X1 U27 ( .A(n119), .B(n146), .Y(n13) );
  MUX2IXL U28 ( .D0(n18), .D1(n52), .S(n148), .Y(n45) );
  AO21X1 U29 ( .B(ps_dat5b[0]), .C(n58), .A(n57), .Y(n59) );
  INVXL U30 ( .A(n103), .Y(k0_det) );
  NAND21XL U31 ( .B(n123), .A(n12), .Y(n124) );
  MUX2BXL U32 ( .D0(n2), .D1(n37), .S(n148), .Y(n14) );
  NAND32XL U33 ( .B(n174), .C(n43), .A(n42), .Y(n56) );
  AND2XL U34 ( .A(prx_fifowdat[5]), .B(prx_fifowdat[7]), .Y(n15) );
  INVX1 U35 ( .A(n41), .Y(n18) );
  NAND31X1 U36 ( .C(n52), .A(n51), .B(n50), .Y(n53) );
  NAND32X1 U37 ( .B(n1), .C(prx_fsm[2]), .A(n170), .Y(n17) );
  NAND31X1 U38 ( .C(bcnt[1]), .A(bcnt[2]), .B(n101), .Y(n104) );
  NAND3XL U39 ( .A(n243), .B(n244), .C(prx_rcvdords[2]), .Y(n224) );
  NAND3XL U40 ( .A(prx_rcvdords[0]), .B(n226), .C(ordsbuf[3]), .Y(n234) );
  INVXL U41 ( .A(prx_rcvdords[1]), .Y(n226) );
  MUX3XL U42 ( .D0(n192), .D1(n191), .D2(n190), .S0(prx_rcvdords[1]), .S1(
        prx_rcvdords[2]), .Y(cs_ords_ena) );
  MUX2XL U43 ( .D0(r_ords_ena[1]), .D1(r_ords_ena[2]), .S(prx_rcvdords[0]), 
        .Y(n191) );
  MUX4XL U44 ( .D0(r_ords_ena[3]), .D1(r_ords_ena[4]), .D2(r_ords_ena[5]), 
        .D3(r_ords_ena[6]), .S0(prx_rcvdords[0]), .S1(prx_rcvdords[1]), .Y(
        n190) );
  INVXL U45 ( .A(prx_rcvdords[2]), .Y(n232) );
  NAND3XL U46 ( .A(n237), .B(n227), .C(prx_rcvdords[1]), .Y(n208) );
  INVXL U47 ( .A(prx_rcvdords[0]), .Y(n193) );
  NAND4XL U48 ( .A(prx_rcvdords[2]), .B(n225), .C(prx_fifowdat[2]), .D(n240), 
        .Y(n200) );
  NAND21X1 U49 ( .B(n248), .A(n92), .Y(n245) );
  INVX1 U50 ( .A(n100), .Y(n92) );
  INVX1 U51 ( .A(n93), .Y(n91) );
  INVX1 U52 ( .A(n81), .Y(n75) );
  INVX1 U53 ( .A(n70), .Y(n72) );
  INVX1 U54 ( .A(n257), .Y(n99) );
  NAND21X1 U55 ( .B(n149), .A(n12), .Y(N153) );
  NOR2X1 U56 ( .A(pid_goidle), .B(n122), .Y(n9) );
  INVX1 U57 ( .A(n143), .Y(n158) );
  INVX1 U58 ( .A(srstz), .Y(n30) );
  INVX1 U59 ( .A(n147), .Y(n133) );
  NAND32X1 U60 ( .B(n131), .C(n30), .A(n150), .Y(N70) );
  INVX1 U61 ( .A(n150), .Y(n152) );
  NOR2X1 U62 ( .A(n88), .B(n11), .Y(n10) );
  OA21X1 U63 ( .B(n247), .C(n223), .A(n248), .Y(n11) );
  INVX1 U64 ( .A(n166), .Y(n168) );
  NAND21X1 U65 ( .B(n195), .A(n13), .Y(n166) );
  INVX1 U66 ( .A(n96), .Y(n69) );
  INVX1 U67 ( .A(N31), .Y(n184) );
  INVX1 U68 ( .A(n88), .Y(n95) );
  NAND21X1 U69 ( .B(n113), .A(n69), .Y(n100) );
  OR2X1 U70 ( .A(n100), .B(n90), .Y(n93) );
  OAI211X1 U71 ( .C(n215), .D(n84), .A(n183), .B(n204), .Y(N33) );
  INVX1 U72 ( .A(n213), .Y(n84) );
  NAND32X1 U73 ( .B(n115), .C(n90), .A(n76), .Y(n81) );
  AO22X1 U74 ( .A(n159), .B(n9), .C(n158), .D(n157), .Y(N276) );
  INVX1 U75 ( .A(n153), .Y(n159) );
  AO21X1 U76 ( .B(n156), .C(n179), .A(n155), .Y(n157) );
  INVX1 U77 ( .A(n154), .Y(n156) );
  OA21X1 U78 ( .B(n141), .C(n140), .A(n158), .Y(N277) );
  OA21X1 U79 ( .B(n139), .C(n140), .A(n158), .Y(N279) );
  INVX1 U80 ( .A(n167), .Y(n117) );
  INVX1 U81 ( .A(n83), .Y(n183) );
  AO21X1 U82 ( .B(n21), .C(n178), .A(prx_setsta[6]), .Y(prx_fiforst) );
  NAND2X1 U83 ( .A(n238), .B(n237), .Y(n70) );
  INVX1 U84 ( .A(n199), .Y(n71) );
  NAND21X1 U85 ( .B(n30), .A(n160), .Y(n122) );
  NOR2X1 U86 ( .A(n122), .B(pid_gobusy), .Y(n12) );
  INVX1 U87 ( .A(n124), .Y(n149) );
  NAND43X1 U88 ( .B(pid_goidle), .C(n30), .D(n117), .A(n21), .Y(n143) );
  NAND32X1 U89 ( .B(n21), .C(n30), .A(n121), .Y(N236) );
  INVXL U90 ( .A(n120), .Y(N251) );
  INVX1 U91 ( .A(n135), .Y(n169) );
  NAND32X1 U92 ( .B(n178), .C(n138), .A(n134), .Y(n155) );
  NAND21X1 U93 ( .B(n178), .A(n111), .Y(n141) );
  AND2X1 U94 ( .A(n133), .B(n132), .Y(N249) );
  INVX1 U95 ( .A(n134), .Y(n139) );
  INVX1 U96 ( .A(n177), .Y(n123) );
  NAND32X1 U97 ( .B(n106), .C(n114), .A(n63), .Y(n103) );
  OAI21BBX1 U98 ( .A(n38), .B(n66), .C(n14), .Y(N96) );
  INVX1 U99 ( .A(n165), .Y(n170) );
  NAND21X1 U100 ( .B(n164), .A(n21), .Y(n165) );
  INVX1 U101 ( .A(n34), .Y(n32) );
  INVX1 U102 ( .A(n182), .Y(prx_cccnt[0]) );
  INVX1 U103 ( .A(n42), .Y(n65) );
  INVX1 U104 ( .A(n64), .Y(n52) );
  NAND32X1 U105 ( .B(n108), .C(n110), .A(n164), .Y(n147) );
  INVX1 U106 ( .A(n146), .Y(n136) );
  OAI221X1 U107 ( .A(n223), .B(n94), .C(n224), .D(n93), .E(n203), .Y(n222) );
  AOI221XL U108 ( .A(n77), .B(n92), .C(n91), .D(n228), .E(n229), .Y(n94) );
  AO21XL U109 ( .B(n169), .C(n21), .A(n168), .Y(prx_crcstart) );
  OAI21AX1 U110 ( .B(n129), .C(n130), .A(n131), .Y(n150) );
  NAND31X1 U111 ( .C(n96), .A(n252), .B(n132), .Y(n88) );
  NAND21X1 U112 ( .B(pff_txreq), .A(n128), .Y(n131) );
  AO21X1 U113 ( .B(N61), .C(n152), .A(n30), .Y(N75) );
  AO21X1 U114 ( .B(N60), .C(n152), .A(n30), .Y(N74) );
  AO21X1 U115 ( .B(N59), .C(n152), .A(n30), .Y(N73) );
  AO21X1 U116 ( .B(N58), .C(n152), .A(n30), .Y(N72) );
  OAI21BBX1 U117 ( .A(n152), .B(n151), .C(srstz), .Y(N71) );
  OAI21AX1 U118 ( .B(n245), .C(n223), .A(n73), .Y(n205) );
  OAI211X1 U119 ( .C(n220), .D(n205), .A(n204), .B(n185), .Y(N31) );
  NAND32X1 U120 ( .B(n82), .C(n83), .A(n217), .Y(N32) );
  INVX1 U121 ( .A(n204), .Y(n82) );
  AO21X1 U122 ( .B(n170), .C(n167), .A(n168), .Y(prx_crcshfi4) );
  AND2XL U123 ( .A(n13), .B(n179), .Y(prx_setsta[2]) );
  INVX1 U124 ( .A(ps_ords_ena), .Y(n179) );
  AND2XL U125 ( .A(ps_ords_ena), .B(n13), .Y(prx_setsta[1]) );
  OAI221X1 U126 ( .A(n216), .B(n97), .C(n96), .D(n98), .E(n207), .Y(n231) );
  AOI32X1 U127 ( .A(n257), .B(n95), .C(n113), .D(n256), .E(n238), .Y(n97) );
  INVX1 U128 ( .A(n221), .Y(n185) );
  NAND43X1 U129 ( .B(n115), .C(n114), .D(prx_fifowdat[5]), .A(n113), .Y(n167)
         );
  INVX1 U130 ( .A(n74), .Y(n76) );
  OAI211X1 U131 ( .C(n224), .D(n81), .A(n200), .B(n80), .Y(n83) );
  AO21X1 U132 ( .B(n79), .C(n78), .A(n239), .Y(n80) );
  INVX1 U133 ( .A(n229), .Y(n78) );
  NAND32X1 U134 ( .B(n169), .C(n138), .A(n137), .Y(n140) );
  AOI32X1 U135 ( .A(n197), .B(ps_ords_ena), .C(n136), .D(n139), .E(n210), .Y(
        n137) );
  AND3X1 U136 ( .A(prx_eoprcvd), .B(pcc_rxgood), .C(n180), .Y(prx_setsta[3])
         );
  AOI21X1 U137 ( .B(n145), .C(n144), .A(n143), .Y(N278) );
  AO21X1 U138 ( .B(ps_ords_ena), .C(n142), .A(n154), .Y(n145) );
  INVX1 U139 ( .A(n195), .Y(n142) );
  INVX1 U140 ( .A(n163), .Y(prx_eoprcvd) );
  NAND32X1 U141 ( .B(n164), .C(n162), .A(n161), .Y(n163) );
  INVX1 U142 ( .A(cs_ords_ena), .Y(n162) );
  INVX1 U143 ( .A(n160), .Y(n161) );
  NAND21X1 U144 ( .B(n146), .A(n197), .Y(n154) );
  INVX1 U145 ( .A(n172), .Y(prx_setsta[6]) );
  NAND32X1 U146 ( .B(n180), .C(n181), .A(prx_eoprcvd), .Y(n172) );
  OAI22AX1 U147 ( .D(N33), .C(n146), .A(n3), .B(n147), .Y(N248) );
  OAI22X1 U148 ( .A(n219), .B(n147), .C(n184), .D(n146), .Y(N246) );
  OAI22AX1 U149 ( .D(N32), .C(n146), .A(n216), .B(n147), .Y(N247) );
  INVX1 U150 ( .A(n212), .Y(n132) );
  AND2X1 U151 ( .A(prx_eoprcvd), .B(n181), .Y(prx_setsta[4]) );
  INVXL U152 ( .A(prx_fifowdat[4]), .Y(n25) );
  NAND43X1 U153 ( .B(n3), .C(n219), .D(prx_rxcode[1]), .A(prx_fifowdat[3]), 
        .Y(n90) );
  BUFXL U154 ( .A(prx_fifowdat[5]), .Y(prx_crcsidat[1]) );
  INVXL U155 ( .A(prx_fifowdat[6]), .Y(n28) );
  NAND21X1 U156 ( .B(n248), .A(n256), .Y(n98) );
  INVX1 U157 ( .A(n224), .Y(n77) );
  OAI211X1 U158 ( .C(n118), .D(n143), .A(n153), .B(n9), .Y(N275) );
  AND4X1 U159 ( .A(n112), .B(n111), .C(n135), .D(n146), .Y(n118) );
  INVX1 U160 ( .A(n155), .Y(n112) );
  OAI211X1 U161 ( .C(n194), .D(n106), .A(srstz), .B(n105), .Y(n121) );
  INVX1 U162 ( .A(pcc_rxgood), .Y(n181) );
  INVX1 U163 ( .A(n106), .Y(n178) );
  NAND21X1 U164 ( .B(n164), .A(n19), .Y(n135) );
  NAND32X1 U165 ( .B(n116), .C(n173), .A(n211), .Y(n153) );
  INVX1 U166 ( .A(pid_gobusy), .Y(n116) );
  INVX1 U167 ( .A(n109), .Y(n138) );
  NAND32X1 U168 ( .B(n108), .C(n141), .A(n110), .Y(n109) );
  INVX1 U169 ( .A(n107), .Y(n111) );
  NAND21X1 U170 ( .B(n133), .A(n144), .Y(n107) );
  NAND32X1 U171 ( .B(n164), .C(n110), .A(n171), .Y(n134) );
  INVX1 U172 ( .A(n194), .Y(n175) );
  AND4XL U173 ( .A(n178), .B(n177), .C(n176), .D(n175), .Y(prx_setsta[0]) );
  INVX1 U174 ( .A(n173), .Y(prx_idle) );
  AND2X1 U175 ( .A(cccnt[3]), .B(cccnt[2]), .Y(n102) );
  INVXL U176 ( .A(n56), .Y(n61) );
  MUX2BX1 U177 ( .D0(n39), .D1(n16), .S(prx_bmc), .Y(n47) );
  NAND4XL U178 ( .A(n148), .B(n66), .C(n43), .D(n44), .Y(n16) );
  INVX1 U179 ( .A(bcnt[0]), .Y(n101) );
  OAI21BBX1 U180 ( .A(r_pshords), .B(N250), .C(n17), .Y(prx_fifopsh) );
  AO21X1 U181 ( .B(cccnt[2]), .C(cccnt[1]), .A(cccnt[5]), .Y(n34) );
  NAND21X1 U182 ( .B(n127), .A(cccnt[4]), .Y(n129) );
  AO21X1 U183 ( .B(shrtrans), .C(n151), .A(n125), .Y(n31) );
  INVX1 U184 ( .A(cccnt[3]), .Y(n127) );
  INVX1 U185 ( .A(n36), .Y(n85) );
  OAI31XL U186 ( .A(n35), .B(cccnt[4]), .C(n34), .D(n33), .Y(n36) );
  AO21X1 U187 ( .B(cccnt[2]), .C(cccnt[0]), .A(cccnt[3]), .Y(n35) );
  AO22X1 U188 ( .A(n32), .B(n31), .C(n129), .D(n126), .Y(n33) );
  INVX1 U189 ( .A(cccnt[0]), .Y(n151) );
  INVX1 U190 ( .A(cccnt[2]), .Y(n125) );
  INVX1 U191 ( .A(cccnt[5]), .Y(n126) );
  NAND32X1 U192 ( .B(cccnt[4]), .C(n130), .A(n127), .Y(n182) );
  NAND42X1 U193 ( .C(n126), .D(n125), .A(cccnt[1]), .B(cccnt[0]), .Y(n130) );
  NAND21X1 U194 ( .B(n66), .A(prx_bmc), .Y(n42) );
  NAND21X1 U195 ( .B(ps_dat5b[2]), .A(ps_dat5b[1]), .Y(n64) );
  AND3X1 U196 ( .A(ps_dat5b[0]), .B(ps_dat5b[2]), .C(n65), .Y(n37) );
  INVX1 U197 ( .A(prx_bmc), .Y(n58) );
  INVX1 U198 ( .A(ps_dat5b[1]), .Y(n66) );
  INVX1 U199 ( .A(ps_dat5b[2]), .Y(n43) );
  INVX1 U200 ( .A(n40), .Y(n48) );
  NAND21X1 U201 ( .B(ps_dat5b[1]), .A(ps_dat5b[2]), .Y(n40) );
  INVX1 U202 ( .A(ps_dat5b[0]), .Y(n44) );
  INVX1 U203 ( .A(shrtrans), .Y(n87) );
  NAND32X1 U204 ( .B(n6), .C(n108), .A(n110), .Y(n106) );
  NAND21X1 U205 ( .B(prx_fsm[2]), .A(prx_fsm[0]), .Y(n108) );
  NAND21X1 U206 ( .B(prx_fsm[3]), .A(n19), .Y(n146) );
  NOR3XL U207 ( .A(n171), .B(n110), .C(prx_fsm[0]), .Y(n19) );
  INVX1 U208 ( .A(prx_fsm[1]), .Y(n110) );
  INVX1 U209 ( .A(prx_fsm[2]), .Y(n171) );
  INVX1 U210 ( .A(prx_fsm[3]), .Y(n164) );
  AOI32X1 U211 ( .A(n236), .B(n237), .C(n69), .D(n10), .E(n216), .Y(n68) );
  MUX2XL U212 ( .D0(N96), .D1(prx_crcsidat[3]), .S(prx_fsm[3]), .Y(
        prx_fifowdat[7]) );
  INVX1 U213 ( .A(n25), .Y(prx_crcsidat[0]) );
  INVX1 U214 ( .A(n67), .Y(prx_crcsidat[3]) );
  AO21X1 U215 ( .B(N62), .C(n152), .A(n30), .Y(N76) );
  INVX1 U216 ( .A(n28), .Y(prx_crcsidat[2]) );
  MUX3X1 U217 ( .D0(n189), .D1(n188), .D2(n187), .S0(N32), .S1(N33), .Y(
        ps_ords_ena) );
  NOR21XL U218 ( .B(r_ords_ena[0]), .A(n184), .Y(n189) );
  MUX2X1 U219 ( .D0(r_ords_ena[1]), .D1(r_ords_ena[2]), .S(N31), .Y(n188) );
  MUX4X1 U220 ( .D0(r_ords_ena[3]), .D1(r_ords_ena[4]), .D2(r_ords_ena[5]), 
        .D3(r_ords_ena[6]), .S0(N31), .S1(N32), .Y(n187) );
  OAI221X1 U221 ( .A(prx_fifowdat[1]), .B(n89), .C(n249), .D(n245), .E(n208), 
        .Y(n218) );
  OA21X1 U222 ( .B(n100), .C(n99), .A(n98), .Y(n262) );
  NOR21XL U223 ( .B(r_ords_ena[0]), .A(n193), .Y(n192) );
  AND2X1 U224 ( .A(n149), .B(prx_bmc), .Y(N156) );
  AND2X1 U225 ( .A(n149), .B(ps_dat5b[2]), .Y(N155) );
  AND2X1 U226 ( .A(n149), .B(ps_dat5b[1]), .Y(N154) );
  INVX1 U227 ( .A(r_rgdcrc), .Y(n180) );
  AO21X1 U228 ( .B(bcnt[0]), .C(bcnt[1]), .A(n121), .Y(n265) );
  NAND21X1 U229 ( .B(n266), .A(bcnt[1]), .Y(n264) );
  NAND21X1 U230 ( .B(n121), .A(bcnt[0]), .Y(n266) );
  NOR2X1 U231 ( .A(bcnt[0]), .B(n121), .Y(n20) );
  NAND21X1 U232 ( .B(shrtrans), .A(n85), .Y(n86) );
  AND3X1 U233 ( .A(pid_goidle), .B(prx_fsm[3]), .C(cs_ords_ena), .Y(
        prx_setsta[5]) );
  NAND43X1 U234 ( .B(prx_fsm[3]), .C(prx_fsm[2]), .D(n110), .A(n210), .Y(n144)
         );
  NAND43X1 U235 ( .B(prx_fsm[1]), .C(prx_fsm[3]), .D(prx_fsm[2]), .A(n210), 
        .Y(n173) );
  NOR21XL U236 ( .B(ps_dat5b[0]), .A(n57), .Y(n55) );
  INVXL U237 ( .A(n57), .Y(n39) );
  NAND32XL U238 ( .B(n66), .C(n43), .A(n174), .Y(n57) );
  AND2XL U239 ( .A(n149), .B(n148), .Y(N157) );
  MUX2IXL U240 ( .D0(ps_dat5b[1]), .D1(n48), .S(n148), .Y(n51) );
  AND3XL U241 ( .A(ps_dat5b[0]), .B(n148), .C(n66), .Y(n60) );
  NAND21X1 U242 ( .B(n49), .A(ps_dat5b[0]), .Y(n50) );
  NAND21X1 U243 ( .B(n268), .A(n62), .Y(n63) );
  INVXL U244 ( .A(n49), .Y(n38) );
  NAND21XL U245 ( .B(n119), .A(n117), .Y(n160) );
  AND3XL U246 ( .A(n119), .B(n177), .C(n173), .Y(n105) );
  MUX2IXL U247 ( .D0(cctrans), .D1(prx_cccnt[0]), .S(n8), .Y(n128) );
  MUX2XL U248 ( .D0(n87), .D1(n86), .S(cctrans), .Y(n196) );
  GEN2XL U249 ( .D(n102), .E(cccnt[4]), .C(cccnt[5]), .B(cctrans), .A(n148), 
        .Y(n177) );
  AOI32XL U250 ( .A(prx_fifowdat[6]), .B(n77), .C(n76), .D(n228), .E(n75), .Y(
        n79) );
  INVXL U251 ( .A(n267), .Y(n115) );
  NAND21XL U252 ( .B(n267), .A(n15), .Y(n96) );
  OAI221XL U253 ( .A(prx_fifowdat[1]), .B(n70), .C(prx_fifowdat[4]), .D(n68), 
        .E(n201), .Y(n221) );
  NAND21XL U254 ( .B(n268), .A(n15), .Y(n74) );
  GEN2XL U255 ( .D(n10), .E(n268), .C(n72), .B(prx_rxcode[1]), .A(n71), .Y(n73) );
  AOI32XL U256 ( .A(n254), .B(n95), .C(n268), .D(n246), .E(n238), .Y(n89) );
  INVXL U257 ( .A(n268), .Y(n113) );
  XOR2XL U258 ( .A(n174), .B(prx_bmc), .Y(n176) );
  GEN2XL U259 ( .D(n263), .E(n66), .C(n65), .B(n64), .A(n174), .Y(n67) );
  NAND21X1 U260 ( .B(n13), .A(n120), .Y(N250) );
  AO21X4 U261 ( .B(n104), .C(n103), .A(n123), .Y(n119) );
  XOR2X1 U262 ( .A(add_83_carry[5]), .B(cccnt[5]), .Y(N62) );
  NOR2X1 U263 ( .A(n30), .B(n196), .Y(n214) );
  NOR2X1 U264 ( .A(n184), .B(n197), .Y(prx_rst[0]) );
  NOR2X1 U265 ( .A(N31), .B(n197), .Y(prx_rst[1]) );
  NOR4XL U266 ( .A(n198), .B(cccnt[2]), .C(cccnt[5]), .D(cccnt[3]), .Y(
        prx_cccnt[1]) );
  NAND3X1 U267 ( .A(cccnt[4]), .B(cccnt[1]), .C(cccnt[0]), .Y(n198) );
  NOR43XL U268 ( .B(n199), .C(n200), .D(n201), .A(n202), .Y(n195) );
  OAI221X1 U269 ( .A(n203), .B(n204), .C(n205), .D(n206), .E(n207), .Y(n202)
         );
  AND2X1 U270 ( .A(n208), .B(n209), .Y(n206) );
  NAND2X1 U271 ( .A(N33), .B(N32), .Y(n197) );
  INVX1 U272 ( .A(n8), .Y(n211) );
  OAI21X1 U273 ( .B(n205), .C(n218), .A(n185), .Y(n217) );
  NAND4X1 U274 ( .A(n183), .B(n213), .C(n215), .D(n222), .Y(n204) );
  NAND3X1 U275 ( .A(n225), .B(n226), .C(n227), .Y(n203) );
  NOR2X1 U276 ( .A(n230), .B(n231), .Y(n215) );
  NOR3XL U277 ( .A(n221), .B(n205), .C(n218), .Y(n213) );
  NAND4X1 U278 ( .A(n219), .B(n3), .C(n232), .D(n233), .Y(n201) );
  NOR3XL U279 ( .A(n223), .B(n234), .C(n235), .Y(n233) );
  NOR3XL U280 ( .A(n235), .B(prx_fifowdat[0]), .C(n234), .Y(n240) );
  INVX1 U281 ( .A(n239), .Y(n225) );
  NAND4X1 U282 ( .A(ordsbuf[7]), .B(ordsbuf[6]), .C(ordsbuf[4]), .D(n241), .Y(
        n239) );
  NOR43XL U283 ( .B(prx_fifowdat[3]), .C(n216), .D(n242), .A(n3), .Y(n229) );
  NOR2X1 U284 ( .A(n219), .B(n224), .Y(n242) );
  OAI21X1 U285 ( .B(n234), .C(n232), .A(r_ordrs4), .Y(n228) );
  NAND3X1 U286 ( .A(n246), .B(n226), .C(n227), .Y(n199) );
  AOI21BX1 U287 ( .C(n230), .B(n231), .A(n218), .Y(n220) );
  NOR43XL U288 ( .B(prx_rcvdords[0]), .C(n232), .D(n250), .A(n251), .Y(n227)
         );
  NOR21XL U289 ( .B(n252), .A(n235), .Y(n250) );
  INVX1 U290 ( .A(n223), .Y(n237) );
  NAND2X1 U291 ( .A(n253), .B(n241), .Y(n223) );
  INVX1 U292 ( .A(ordsbuf[5]), .Y(n241) );
  OAI21X1 U293 ( .B(n247), .C(n249), .A(n248), .Y(n254) );
  NAND4X1 U294 ( .A(n255), .B(n246), .C(n193), .D(n219), .Y(n207) );
  INVX1 U295 ( .A(n249), .Y(n246) );
  NAND2X1 U296 ( .A(ordsbuf[5]), .B(n253), .Y(n249) );
  NOR32XL U297 ( .B(ordsbuf[4]), .C(ordsbuf[7]), .A(ordsbuf[6]), .Y(n253) );
  NOR32XL U298 ( .B(prx_fifowdat[3]), .C(n252), .A(n248), .Y(n238) );
  NOR2X1 U299 ( .A(n219), .B(n269), .Y(n252) );
  OAI211X1 U300 ( .C(n245), .D(n258), .A(n259), .B(n209), .Y(n230) );
  NAND4X1 U301 ( .A(n256), .B(n255), .C(prx_fifowdat[0]), .D(n193), .Y(n209)
         );
  NOR32XL U302 ( .B(prx_rcvdords[1]), .C(n260), .A(n232), .Y(n255) );
  NOR3XL U303 ( .A(n235), .B(prx_fifowdat[2]), .C(n251), .Y(n260) );
  INVX1 U304 ( .A(ordsbuf[3]), .Y(n251) );
  NAND32X1 U305 ( .B(r_exist1st), .C(n216), .A(prx_fifowdat[3]), .Y(n235) );
  INVX1 U306 ( .A(prx_fifowdat[1]), .Y(n216) );
  NAND4X1 U307 ( .A(prx_fifowdat[2]), .B(prx_fifowdat[1]), .C(n261), .D(
        prx_fifowdat[3]), .Y(n259) );
  INVX1 U308 ( .A(n212), .Y(prx_fifowdat[3]) );
  MUX2IX1 U309 ( .D0(prx_rxcode[4]), .D1(prx_rxcode[3]), .S(prx_fsm[3]), .Y(
        n212) );
  NOR2X1 U310 ( .A(prx_fifowdat[0]), .B(n262), .Y(n261) );
  OAI21X1 U311 ( .B(n247), .C(n258), .A(n248), .Y(n257) );
  AOI21X1 U312 ( .B(n232), .C(n243), .A(n244), .Y(n247) );
  INVX1 U313 ( .A(n256), .Y(n258) );
  NOR43XL U314 ( .B(ordsbuf[6]), .C(ordsbuf[7]), .D(ordsbuf[5]), .A(ordsbuf[4]), .Y(n256) );
  INVX1 U315 ( .A(n248), .Y(n236) );
  NAND3X1 U316 ( .A(n232), .B(n244), .C(n243), .Y(n248) );
  INVX1 U317 ( .A(n234), .Y(n243) );
  INVX1 U318 ( .A(r_ordrs4), .Y(n244) );
  NAND2X1 U319 ( .A(prx_bmc), .B(ps_dat5b[2]), .Y(n263) );
  INVX1 U320 ( .A(prx_fifowdat[0]), .Y(n219) );
  MUX2IX1 U321 ( .D0(n264), .D1(n265), .S(bcnt[2]), .Y(N239) );
  MUX2AXL U322 ( .D0(n266), .D1(n20), .S(bcnt[1]), .Y(N238) );
  NOR2X1 U323 ( .A(bcnt[2]), .B(bcnt[1]), .Y(n194) );
  INVX1 U324 ( .A(prx_fsm[0]), .Y(n210) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyrx_a0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyrx_a0_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyrx_a0_3 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyrx_a0_4 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyrx_a0_5 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyrx_a0_6 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyrx_a0_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module phyrx_adp ( clk, srstz, gohi, golo, gobusy, goidle, i_ccidle, k0_det, 
        r_adprx_en, r_adp2nd, adp_val, d_cc, cctrans );
  output [5:0] adp_val;
  input clk, srstz, gohi, golo, gobusy, goidle, i_ccidle, k0_det, r_adprx_en,
         r_adp2nd;
  output d_cc, cctrans;
  wire   N49, N50, N51, N52, N53, N54, N55, N70, N71, N72, N73, N74, N97, N98,
         N99, N100, N101, N102, N103, N104, N106, N107, N108, N109, N110, N111,
         N112, N130, N131, N132, N133, N134, N135, N136, N137, N138, N139,
         N140, N141, N142, N143, N144, N145, N169, N170, N171, N172, N173,
         net10687, net10693, net10698, net10703, n115, n1, n2, n3, n4, n5, n6,
         n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112,
         SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2,
         SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4,
         SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6,
         SYNOPSYS_UNCONNECTED_7;
  wire   [7:0] dcnt_h;
  wire   [5:0] adp_v0;
  wire   [3:0] dcnt_n;
  wire   [5:0] dcnt_e;

  SNPS_CLOCK_GATE_HIGH_phyrx_adp_0 clk_gate_adp_n_reg ( .CLK(clk), .EN(N49), 
        .ENCLK(net10687), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_phyrx_adp_3 clk_gate_dcnt_e_reg ( .CLK(clk), .EN(N130), 
        .ENCLK(net10693), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_phyrx_adp_2 clk_gate_dcnt_h_reg ( .CLK(clk), .EN(N137), 
        .ENCLK(net10698), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_phyrx_adp_1 clk_gate_dcnt_n_reg ( .CLK(clk), .EN(N169), 
        .ENCLK(net10703), .TE(1'b0) );
  phyrx_adp_DW01_inc_0 add_385 ( .A({n2, dcnt_h[6:0]}), .SUM({N104, N103, N102, 
        N101, N100, N99, N98, N97}) );
  phyrx_adp_DW_div_tc_6 div_338 ( .a({dcnt_h[7], n2, dcnt_h[6:0]}), .b({1'b0, 
        1'b1, 1'b1, 1'b0}), .quotient({SYNOPSYS_UNCONNECTED_1, 
        SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3, adp_v0}), .remainder({
        SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6, 
        SYNOPSYS_UNCONNECTED_7}), .divide_by_0() );
  DFFQX1 dcnt_h_reg_6_ ( .D(N144), .C(net10698), .Q(dcnt_h[6]) );
  DFFQX1 dcnt_h_reg_4_ ( .D(N142), .C(net10698), .Q(dcnt_h[4]) );
  DFFQX1 dcnt_h_reg_5_ ( .D(N143), .C(net10698), .Q(dcnt_h[5]) );
  DFFQX1 dcnt_h_reg_1_ ( .D(N139), .C(net10698), .Q(dcnt_h[1]) );
  DFFQX1 dcnt_h_reg_2_ ( .D(N140), .C(net10698), .Q(dcnt_h[2]) );
  DFFQX1 dcnt_h_reg_3_ ( .D(N141), .C(net10698), .Q(dcnt_h[3]) );
  DFFQX1 dcnt_h_reg_0_ ( .D(N138), .C(net10698), .Q(dcnt_h[0]) );
  DFFQX1 dcnt_h_reg_7_ ( .D(N145), .C(net10698), .Q(dcnt_h[7]) );
  DFFQX1 adp_n_reg_5_ ( .D(N55), .C(net10687), .Q(adp_val[5]) );
  DFFQX1 dcnt_n_reg_2_ ( .D(N172), .C(net10703), .Q(dcnt_n[2]) );
  DFFQX1 dcnt_n_reg_1_ ( .D(N171), .C(net10703), .Q(dcnt_n[1]) );
  DFFQX1 adp_n_reg_4_ ( .D(N54), .C(net10687), .Q(adp_val[4]) );
  DFFQX1 adp_n_reg_2_ ( .D(N52), .C(net10687), .Q(adp_val[2]) );
  DFFQX1 dcnt_e_reg_0_ ( .D(N131), .C(net10693), .Q(dcnt_e[0]) );
  DFFQX1 cs_d_cc_reg ( .D(n115), .C(clk), .Q(d_cc) );
  DFFQX1 adp_n_reg_3_ ( .D(N53), .C(net10687), .Q(adp_val[3]) );
  DFFQX1 dcnt_n_reg_3_ ( .D(N173), .C(net10703), .Q(dcnt_n[3]) );
  DFFQX1 dcnt_n_reg_0_ ( .D(N170), .C(net10703), .Q(dcnt_n[0]) );
  DFFQX1 adp_n_reg_1_ ( .D(N51), .C(net10687), .Q(adp_val[1]) );
  DFFQX1 adp_n_reg_0_ ( .D(N50), .C(net10687), .Q(adp_val[0]) );
  DFFQX1 dcnt_e_reg_3_ ( .D(N134), .C(net10693), .Q(dcnt_e[3]) );
  DFFQX1 dcnt_e_reg_2_ ( .D(N133), .C(net10693), .Q(dcnt_e[2]) );
  DFFQX1 dcnt_e_reg_5_ ( .D(N136), .C(net10693), .Q(dcnt_e[5]) );
  DFFQX1 dcnt_e_reg_1_ ( .D(N132), .C(net10693), .Q(dcnt_e[1]) );
  DFFQX1 dcnt_e_reg_4_ ( .D(N135), .C(net10693), .Q(dcnt_e[4]) );
  INVX1 U3 ( .A(golo), .Y(n12) );
  NOR21XL U4 ( .B(n89), .A(n36), .Y(n37) );
  AND2X1 U5 ( .A(dcnt_e[4]), .B(dcnt_e[2]), .Y(n1) );
  BUFX3 U6 ( .A(dcnt_h[7]), .Y(n2) );
  MUX2IX2 U7 ( .D0(n12), .D1(n13), .S(n58), .Y(n6) );
  INVX1 U8 ( .A(n3), .Y(n65) );
  NAND21X1 U9 ( .B(n13), .A(adp_val[4]), .Y(n15) );
  XNOR2XL U10 ( .A(dcnt_e[4]), .B(dcnt_e[5]), .Y(n52) );
  OR3XL U11 ( .A(dcnt_e[3]), .B(dcnt_e[2]), .C(dcnt_e[1]), .Y(n29) );
  NAND3XL U12 ( .A(n39), .B(n35), .C(n37), .Y(n63) );
  NAND43XL U13 ( .B(n89), .C(n11), .D(n40), .A(n39), .Y(n62) );
  NAND21XL U14 ( .B(n64), .A(n4), .Y(n3) );
  NAND4X1 U15 ( .A(dcnt_e[0]), .B(dcnt_e[1]), .C(dcnt_e[3]), .D(n1), .Y(n4) );
  MUX2IX1 U16 ( .D0(n15), .D1(n14), .S(d_cc), .Y(n26) );
  NOR31X1 U17 ( .C(n22), .A(adp_val[0]), .B(n21), .Y(n23) );
  AOI22XL U18 ( .A(n92), .B(dcnt_e[0]), .C(n91), .D(dcnt_e[5]), .Y(n48) );
  OR2XL U19 ( .A(dcnt_e[3]), .B(n51), .Y(n45) );
  INVXL U20 ( .A(n52), .Y(n27) );
  OR2XL U21 ( .A(dcnt_e[4]), .B(n70), .Y(n71) );
  OAI21BBXL U22 ( .A(n68), .B(dcnt_e[2]), .C(n69), .Y(N71) );
  OAI21BBXL U23 ( .A(dcnt_e[0]), .B(dcnt_e[1]), .C(n68), .Y(N70) );
  NAND2XL U24 ( .A(dcnt_e[0]), .B(n53), .Y(n44) );
  OR2XL U25 ( .A(dcnt_e[5]), .B(n30), .Y(n32) );
  INVXL U26 ( .A(dcnt_e[4]), .Y(n91) );
  INVXL U27 ( .A(dcnt_e[0]), .Y(n46) );
  OR2XL U28 ( .A(n69), .B(dcnt_e[3]), .Y(n70) );
  OR2XL U29 ( .A(dcnt_e[1]), .B(dcnt_e[0]), .Y(n68) );
  OR2XL U30 ( .A(n68), .B(dcnt_e[2]), .Y(n69) );
  INVX1 U31 ( .A(n11), .Y(n10) );
  INVX1 U32 ( .A(srstz), .Y(n11) );
  AO21X1 U33 ( .B(n47), .C(n43), .A(k0_det), .Y(n51) );
  NAND43X1 U34 ( .B(n41), .C(n55), .D(n40), .A(n10), .Y(N169) );
  INVX1 U35 ( .A(n63), .Y(n41) );
  INVX1 U36 ( .A(n62), .Y(n55) );
  INVX1 U37 ( .A(gohi), .Y(n13) );
  NOR21XL U38 ( .B(n35), .A(n38), .Y(n24) );
  NOR21XL U39 ( .B(n56), .A(n79), .Y(N53) );
  NOR21XL U40 ( .B(n56), .A(n80), .Y(N52) );
  NOR21XL U41 ( .B(n56), .A(n81), .Y(N51) );
  NOR21XL U42 ( .B(n56), .A(n82), .Y(N50) );
  NOR21XL U43 ( .B(n56), .A(n78), .Y(N54) );
  INVX1 U44 ( .A(n57), .Y(n60) );
  NAND32X1 U45 ( .B(n90), .C(n59), .A(n58), .Y(n57) );
  NOR3XL U46 ( .A(n59), .B(n58), .C(n90), .Y(n5) );
  NAND42X1 U47 ( .C(n90), .D(n51), .A(n50), .B(n59), .Y(N137) );
  NAND31X1 U48 ( .C(n44), .A(n52), .B(n47), .Y(n50) );
  AO21X1 U49 ( .B(n9), .C(n7), .A(n34), .Y(n112) );
  INVX1 U50 ( .A(n31), .Y(n67) );
  NAND32X1 U51 ( .B(n34), .C(n7), .A(n9), .Y(n31) );
  INVX1 U52 ( .A(n42), .Y(n47) );
  NAND21X1 U53 ( .B(n56), .A(n10), .Y(N49) );
  NOR21XL U54 ( .B(n55), .A(n87), .Y(N172) );
  OR2X1 U55 ( .A(n91), .B(n44), .Y(n30) );
  INVX1 U56 ( .A(n29), .Y(n53) );
  INVX1 U57 ( .A(n32), .Y(n43) );
  INVX1 U58 ( .A(n38), .Y(n40) );
  NAND21X1 U59 ( .B(n26), .A(n25), .Y(n66) );
  MUX2IX1 U60 ( .D0(n6), .D1(n24), .S(n39), .Y(n25) );
  NAND21XL U61 ( .B(adp_val[4]), .A(golo), .Y(n14) );
  NOR21XL U62 ( .B(n64), .A(n23), .Y(n39) );
  NAND21X1 U63 ( .B(adp_val[3]), .A(n20), .Y(n21) );
  NAND43X1 U64 ( .B(n19), .C(n18), .D(n17), .A(n16), .Y(n38) );
  XOR2X1 U65 ( .A(n22), .B(dcnt_n[2]), .Y(n16) );
  XOR2X1 U66 ( .A(dcnt_n[1]), .B(adp_val[1]), .Y(n19) );
  XOR2X1 U67 ( .A(dcnt_n[3]), .B(adp_val[3]), .Y(n17) );
  OAI31XL U68 ( .A(dcnt_e[0]), .B(dcnt_e[4]), .C(n29), .D(n52), .Y(n64) );
  XOR2X1 U69 ( .A(adp_val[0]), .B(dcnt_n[0]), .Y(n18) );
  XOR2X1 U70 ( .A(n58), .B(adp_val[4]), .Y(n35) );
  INVX1 U71 ( .A(d_cc), .Y(n58) );
  INVX1 U72 ( .A(adp_val[1]), .Y(n20) );
  INVX1 U73 ( .A(adp_val[2]), .Y(n22) );
  AOI32X1 U74 ( .A(n95), .B(n33), .C(n43), .D(N72), .E(n67), .Y(n94) );
  INVX1 U75 ( .A(n34), .Y(n33) );
  NAND21X1 U76 ( .B(n49), .A(n48), .Y(n59) );
  GEN2XL U77 ( .D(n47), .E(n52), .C(n46), .B(n53), .A(n45), .Y(n49) );
  AO22X1 U78 ( .A(N111), .B(n60), .C(N103), .D(n5), .Y(N144) );
  AO22X1 U79 ( .A(N110), .B(n60), .C(N102), .D(n5), .Y(N143) );
  AO22X1 U80 ( .A(N109), .B(n60), .C(N101), .D(n5), .Y(N142) );
  AO22X1 U81 ( .A(N108), .B(n60), .C(N100), .D(n5), .Y(N141) );
  AO22X1 U82 ( .A(N107), .B(n60), .C(N99), .D(n5), .Y(N140) );
  AO22X1 U83 ( .A(N106), .B(n60), .C(N98), .D(n5), .Y(N139) );
  AO22X1 U84 ( .A(N112), .B(n60), .C(N104), .D(n5), .Y(N145) );
  AO22AXL U85 ( .A(N97), .B(n5), .C(n60), .D(dcnt_h[0]), .Y(N138) );
  AO21X1 U86 ( .B(r_adprx_en), .C(k0_det), .A(n42), .Y(n34) );
  NAND21X1 U87 ( .B(i_ccidle), .A(n28), .Y(n42) );
  INVX1 U88 ( .A(n54), .Y(n56) );
  AND2X1 U89 ( .A(n61), .B(n10), .Y(n115) );
  NOR21XL U90 ( .B(n56), .A(dcnt_e[5]), .Y(N55) );
  OAI22X1 U91 ( .A(n11), .B(n63), .C(dcnt_n[0]), .D(n62), .Y(N170) );
  NOR21XL U92 ( .B(n55), .A(n83), .Y(N173) );
  NOR21XL U93 ( .B(n55), .A(n88), .Y(N171) );
  NOR4XL U94 ( .A(dcnt_e[2]), .B(dcnt_e[1]), .C(dcnt_e[0]), .D(n8), .Y(n7) );
  OR3XL U95 ( .A(dcnt_e[3]), .B(dcnt_e[5]), .C(dcnt_e[4]), .Y(n8) );
  OA21X1 U96 ( .B(r_adp2nd), .C(n30), .A(n32), .Y(n9) );
  XOR2XL U97 ( .A(n66), .B(d_cc), .Y(n61) );
  NOR21X2 U98 ( .B(n66), .A(n65), .Y(cctrans) );
  MUX2IXL U99 ( .D0(gohi), .D1(golo), .S(adp_val[4]), .Y(n36) );
  NAND5XL U100 ( .A(n10), .B(dcnt_e[0]), .C(n53), .D(n52), .E(n6), .Y(n54) );
  MUX2XL U101 ( .D0(n6), .D1(n66), .S(n27), .Y(n28) );
  OAI21BBX1 U102 ( .A(n69), .B(dcnt_e[3]), .C(n70), .Y(N72) );
  XNOR2XL U103 ( .A(n70), .B(dcnt_e[4]), .Y(N73) );
  XNOR2XL U104 ( .A(dcnt_e[5]), .B(n71), .Y(N74) );
  OR2X1 U105 ( .A(dcnt_h[1]), .B(dcnt_h[0]), .Y(n72) );
  OAI21BBX1 U106 ( .A(dcnt_h[0]), .B(dcnt_h[1]), .C(n72), .Y(N106) );
  OR2X1 U107 ( .A(n72), .B(dcnt_h[2]), .Y(n73) );
  OAI21BBX1 U108 ( .A(n72), .B(dcnt_h[2]), .C(n73), .Y(N107) );
  OR2X1 U109 ( .A(n73), .B(dcnt_h[3]), .Y(n74) );
  OAI21BBX1 U110 ( .A(n73), .B(dcnt_h[3]), .C(n74), .Y(N108) );
  OR2X1 U111 ( .A(n74), .B(dcnt_h[4]), .Y(n75) );
  OAI21BBX1 U112 ( .A(n74), .B(dcnt_h[4]), .C(n75), .Y(N109) );
  OR2X1 U113 ( .A(n75), .B(dcnt_h[5]), .Y(n76) );
  OAI21BBX1 U114 ( .A(n75), .B(dcnt_h[5]), .C(n76), .Y(N110) );
  XNOR2XL U115 ( .A(n76), .B(dcnt_h[6]), .Y(N111) );
  OR2X1 U116 ( .A(dcnt_h[6]), .B(n76), .Y(n77) );
  XNOR2XL U117 ( .A(n2), .B(n77), .Y(N112) );
  XNOR2XL U118 ( .A(dcnt_n[3]), .B(n84), .Y(n83) );
  NOR2X1 U119 ( .A(n85), .B(n86), .Y(n84) );
  XNOR2XL U120 ( .A(n86), .B(n85), .Y(n87) );
  INVX1 U121 ( .A(dcnt_n[2]), .Y(n85) );
  NAND2X1 U122 ( .A(dcnt_n[1]), .B(dcnt_n[0]), .Y(n86) );
  XNOR2XL U123 ( .A(dcnt_n[1]), .B(dcnt_n[0]), .Y(n88) );
  NOR4XL U124 ( .A(dcnt_n[0]), .B(dcnt_n[1]), .C(dcnt_n[2]), .D(dcnt_n[3]), 
        .Y(n89) );
  AND2X1 U125 ( .A(dcnt_e[1]), .B(dcnt_e[2]), .Y(n92) );
  OAI21BBX1 U126 ( .A(N74), .B(n67), .C(n93), .Y(N136) );
  OAI21BBX1 U127 ( .A(N73), .B(n67), .C(n93), .Y(N135) );
  NAND2X1 U128 ( .A(n94), .B(n93), .Y(N134) );
  OAI211X1 U129 ( .C(n82), .D(n81), .A(n79), .B(n80), .Y(n95) );
  XOR2X1 U130 ( .A(n96), .B(n97), .Y(n80) );
  NOR2X1 U131 ( .A(n98), .B(n78), .Y(n97) );
  XOR2X1 U132 ( .A(n99), .B(n100), .Y(n79) );
  AOI21X1 U133 ( .B(adp_v0[3]), .C(n101), .A(n102), .Y(n100) );
  AOI21X1 U134 ( .B(n98), .C(n96), .A(n78), .Y(n99) );
  OAI21X1 U135 ( .B(adp_v0[2]), .C(n102), .A(n101), .Y(n96) );
  INVX1 U136 ( .A(n103), .Y(n98) );
  NAND2X1 U137 ( .A(n104), .B(n103), .Y(n81) );
  NAND2X1 U138 ( .A(n82), .B(n105), .Y(n103) );
  MUX2IX1 U139 ( .D0(n106), .D1(n78), .S(n105), .Y(n104) );
  OAI21X1 U140 ( .B(adp_v0[1]), .C(n102), .A(n101), .Y(n105) );
  NOR2X1 U141 ( .A(n82), .B(n78), .Y(n106) );
  AOI21BBXL U142 ( .B(n102), .C(n107), .A(n108), .Y(n78) );
  NOR3XL U143 ( .A(adp_v0[0]), .B(n102), .C(n108), .Y(n82) );
  INVX1 U144 ( .A(n101), .Y(n108) );
  OAI21X1 U145 ( .B(n109), .C(n107), .A(adp_v0[5]), .Y(n101) );
  NOR3XL U146 ( .A(adp_v0[1]), .B(adp_v0[3]), .C(adp_v0[2]), .Y(n109) );
  NOR2X1 U147 ( .A(n107), .B(adp_v0[5]), .Y(n102) );
  INVX1 U148 ( .A(adp_v0[4]), .Y(n107) );
  OAI21BBX1 U149 ( .A(N71), .B(n67), .C(n93), .Y(N133) );
  OAI21BBX1 U150 ( .A(N70), .B(n67), .C(n93), .Y(N132) );
  OAI21BBX1 U151 ( .A(n46), .B(n67), .C(n93), .Y(N131) );
  AOI21X1 U152 ( .B(n110), .C(n67), .A(n90), .Y(n93) );
  INVX1 U153 ( .A(n111), .Y(n90) );
  OAI2B11X1 U154 ( .D(k0_det), .C(n110), .A(n112), .B(n111), .Y(N130) );
  NOR3XL U155 ( .A(goidle), .B(gobusy), .C(n11), .Y(n111) );
  INVX1 U156 ( .A(r_adprx_en), .Y(n110) );
endmodule


module phyrx_adp_DW_div_tc_6 ( a, b, quotient, remainder, divide_by_0 );
  input [8:0] a;
  input [3:0] b;
  output [8:0] quotient;
  output [3:0] remainder;
  output divide_by_0;
  wire   u_div_SumTmp_1__0_, u_div_SumTmp_1__2_, u_div_SumTmp_2__0_,
         u_div_SumTmp_3__0_, u_div_SumTmp_4__0_, u_div_SumTmp_5__0_,
         u_div_CryTmp_0__2_, u_div_CryTmp_0__3_, u_div_CryTmp_0__4_,
         u_div_CryTmp_1__2_, u_div_CryTmp_1__4_, u_div_CryTmp_2__4_,
         u_div_CryTmp_3__4_, u_div_CryTmp_4__4_, u_div_CryTmp_5__4_,
         u_div_PartRem_1__2_, u_div_PartRem_1__3_, u_div_PartRem_2__2_,
         u_div_PartRem_2__3_, u_div_PartRem_3__2_, u_div_PartRem_3__3_,
         u_div_PartRem_4__2_, u_div_PartRem_4__3_, u_div_PartRem_5__2_,
         u_div_PartRem_5__3_, u_div_PartRem_7__0_, u_div_PartRem_7__1_, n1, n2,
         n3, n4, n5, n6, n7, n8, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22;
  wire   [5:1] u_div_QIncCry;
  wire   [5:0] u_div_QInv;
  wire   [6:1] u_div_AIncCry;
  wire   [6:0] u_div_AInv;

  HAD1X1 u_div_u_ha_AInc_6 ( .A(u_div_AInv[6]), .B(u_div_AIncCry[6]), .CO(
        u_div_PartRem_7__1_), .SO(u_div_PartRem_7__0_) );
  HAD1X1 u_div_u_ha_AInc_5 ( .A(u_div_AInv[5]), .B(u_div_AIncCry[5]), .CO(
        u_div_AIncCry[6]), .SO(u_div_SumTmp_5__0_) );
  HAD1X1 u_div_u_ha_AInc_4 ( .A(u_div_AInv[4]), .B(u_div_AIncCry[4]), .CO(
        u_div_AIncCry[5]), .SO(u_div_SumTmp_4__0_) );
  HAD1X1 u_div_u_ha_AInc_3 ( .A(u_div_AInv[3]), .B(u_div_AIncCry[3]), .CO(
        u_div_AIncCry[4]), .SO(u_div_SumTmp_3__0_) );
  HAD1X1 u_div_u_ha_AInc_2 ( .A(u_div_AInv[2]), .B(u_div_AIncCry[2]), .CO(
        u_div_AIncCry[3]), .SO(u_div_SumTmp_2__0_) );
  HAD1X1 u_div_u_ha_AInc_1 ( .A(u_div_AInv[1]), .B(u_div_AIncCry[1]), .CO(
        u_div_AIncCry[2]), .SO(u_div_SumTmp_1__0_) );
  HAD1X1 u_div_u_ha_QInc_4 ( .A(u_div_QInv[4]), .B(u_div_QIncCry[4]), .CO(
        u_div_QIncCry[5]), .SO(quotient[4]) );
  HAD1X1 u_div_u_ha_QInc_3 ( .A(u_div_QInv[3]), .B(u_div_QIncCry[3]), .CO(
        u_div_QIncCry[4]), .SO(quotient[3]) );
  HAD1X1 u_div_u_ha_QInc_2 ( .A(u_div_QInv[2]), .B(u_div_QIncCry[2]), .CO(
        u_div_QIncCry[3]), .SO(quotient[2]) );
  HAD1X1 u_div_u_ha_QInc_1 ( .A(u_div_QInv[1]), .B(u_div_QIncCry[1]), .CO(
        u_div_QIncCry[2]), .SO(quotient[1]) );
  HAD1X1 u_div_u_ha_QInc_0 ( .A(u_div_QInv[0]), .B(a[7]), .CO(u_div_QIncCry[1]), .SO(quotient[0]) );
  AND2X1 u_div_u_ha_AInc_0 ( .A(u_div_AInv[0]), .B(a[8]), .Y(u_div_AIncCry[1])
         );
  XOR2X1 u_div_u_ha_QInc_5 ( .A(u_div_QInv[5]), .B(u_div_QIncCry[5]), .Y(
        quotient[5]) );
  NAND2X1 U1 ( .A(u_div_PartRem_4__2_), .B(n11), .Y(n1) );
  NAND2X1 U2 ( .A(u_div_PartRem_3__2_), .B(n12), .Y(n2) );
  NAND2X1 U3 ( .A(u_div_PartRem_5__2_), .B(n10), .Y(n3) );
  NAND2X1 U4 ( .A(u_div_PartRem_2__2_), .B(u_div_CryTmp_1__2_), .Y(n4) );
  XNOR2XL U5 ( .A(n10), .B(u_div_PartRem_5__2_), .Y(n5) );
  XNOR2XL U6 ( .A(n11), .B(u_div_PartRem_4__2_), .Y(n6) );
  XNOR2XL U7 ( .A(n12), .B(u_div_PartRem_3__2_), .Y(n7) );
  XNOR2XL U8 ( .A(u_div_PartRem_7__0_), .B(u_div_PartRem_7__1_), .Y(n8) );
  NAND21X1 U9 ( .B(u_div_PartRem_4__3_), .A(n1), .Y(u_div_CryTmp_3__4_) );
  MUX2IX1 U10 ( .D0(n17), .D1(n5), .S(u_div_CryTmp_4__4_), .Y(
        u_div_PartRem_4__3_) );
  NAND21X1 U11 ( .B(u_div_PartRem_3__3_), .A(n2), .Y(u_div_CryTmp_2__4_) );
  MUX2IX1 U12 ( .D0(n18), .D1(n6), .S(u_div_CryTmp_3__4_), .Y(
        u_div_PartRem_3__3_) );
  NAND21X1 U13 ( .B(u_div_PartRem_2__3_), .A(n4), .Y(u_div_CryTmp_1__4_) );
  MUX2IX1 U14 ( .D0(n19), .D1(n7), .S(u_div_CryTmp_2__4_), .Y(
        u_div_PartRem_2__3_) );
  INVX1 U15 ( .A(n17), .Y(u_div_PartRem_5__2_) );
  INVX1 U16 ( .A(n18), .Y(u_div_PartRem_4__2_) );
  INVX1 U17 ( .A(n19), .Y(u_div_PartRem_3__2_) );
  INVX1 U18 ( .A(n20), .Y(u_div_PartRem_2__2_) );
  MUX2AXL U19 ( .D0(n20), .D1(u_div_SumTmp_1__2_), .S(u_div_CryTmp_1__4_), .Y(
        u_div_PartRem_1__3_) );
  XOR2X1 U20 ( .A(u_div_CryTmp_1__2_), .B(u_div_PartRem_2__2_), .Y(
        u_div_SumTmp_1__2_) );
  AND2X1 U21 ( .A(u_div_PartRem_7__1_), .B(u_div_PartRem_7__0_), .Y(
        u_div_CryTmp_5__4_) );
  MUX2AXL U22 ( .D0(u_div_PartRem_7__0_), .D1(u_div_PartRem_7__0_), .S(
        u_div_CryTmp_5__4_), .Y(n17) );
  MUX2AXL U23 ( .D0(n10), .D1(n10), .S(u_div_CryTmp_4__4_), .Y(n18) );
  MUX2AXL U24 ( .D0(n12), .D1(n12), .S(u_div_CryTmp_2__4_), .Y(n20) );
  MUX2AXL U25 ( .D0(n11), .D1(n11), .S(u_div_CryTmp_3__4_), .Y(n19) );
  MUX2AXL U26 ( .D0(n21), .D1(n21), .S(u_div_CryTmp_1__4_), .Y(
        u_div_PartRem_1__2_) );
  INVX1 U27 ( .A(n21), .Y(u_div_CryTmp_1__2_) );
  INVX1 U28 ( .A(u_div_CryTmp_0__3_), .Y(n13) );
  NOR21XL U29 ( .B(u_div_CryTmp_0__2_), .A(n14), .Y(u_div_CryTmp_0__3_) );
  INVX1 U30 ( .A(u_div_PartRem_1__2_), .Y(n14) );
  MUX2IX1 U31 ( .D0(n22), .D1(n22), .S(u_div_CryTmp_1__4_), .Y(
        u_div_CryTmp_0__2_) );
  NAND21X1 U32 ( .B(u_div_PartRem_5__3_), .A(n3), .Y(u_div_CryTmp_4__4_) );
  MUX2IX1 U33 ( .D0(n16), .D1(n8), .S(u_div_CryTmp_5__4_), .Y(
        u_div_PartRem_5__3_) );
  MUX2IX1 U34 ( .D0(u_div_SumTmp_2__0_), .D1(u_div_SumTmp_2__0_), .S(
        u_div_CryTmp_2__4_), .Y(n21) );
  MUX2X1 U35 ( .D0(u_div_SumTmp_5__0_), .D1(u_div_SumTmp_5__0_), .S(
        u_div_CryTmp_5__4_), .Y(n10) );
  XNOR2XL U36 ( .A(a[7]), .B(n15), .Y(u_div_QInv[5]) );
  INVX1 U37 ( .A(u_div_CryTmp_5__4_), .Y(n15) );
  MUX2X1 U38 ( .D0(u_div_SumTmp_4__0_), .D1(u_div_SumTmp_4__0_), .S(
        u_div_CryTmp_4__4_), .Y(n11) );
  MUX2X1 U39 ( .D0(u_div_SumTmp_3__0_), .D1(u_div_SumTmp_3__0_), .S(
        u_div_CryTmp_3__4_), .Y(n12) );
  INVX1 U40 ( .A(u_div_PartRem_7__1_), .Y(n16) );
  XOR2X1 U41 ( .A(a[7]), .B(u_div_CryTmp_4__4_), .Y(u_div_QInv[4]) );
  XOR2X1 U42 ( .A(a[7]), .B(u_div_CryTmp_0__4_), .Y(u_div_QInv[0]) );
  NAND21X1 U43 ( .B(u_div_PartRem_1__3_), .A(n13), .Y(u_div_CryTmp_0__4_) );
  XOR2X1 U44 ( .A(a[7]), .B(u_div_CryTmp_1__4_), .Y(u_div_QInv[1]) );
  XOR2X1 U45 ( .A(a[7]), .B(u_div_CryTmp_2__4_), .Y(u_div_QInv[2]) );
  XOR2X1 U46 ( .A(a[7]), .B(u_div_CryTmp_3__4_), .Y(u_div_QInv[3]) );
  INVX1 U47 ( .A(u_div_SumTmp_1__0_), .Y(n22) );
  XOR2X1 U48 ( .A(a[8]), .B(a[6]), .Y(u_div_AInv[6]) );
  XOR2X1 U49 ( .A(a[8]), .B(a[1]), .Y(u_div_AInv[1]) );
  XOR2X1 U50 ( .A(a[8]), .B(a[0]), .Y(u_div_AInv[0]) );
  XOR2X1 U51 ( .A(a[8]), .B(a[2]), .Y(u_div_AInv[2]) );
  XOR2X1 U52 ( .A(a[8]), .B(a[3]), .Y(u_div_AInv[3]) );
  XOR2X1 U53 ( .A(a[8]), .B(a[4]), .Y(u_div_AInv[4]) );
  XOR2X1 U54 ( .A(a[8]), .B(a[5]), .Y(u_div_AInv[5]) );
endmodule


module phyrx_adp_DW01_inc_0 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  XOR2X1 U1 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyrx_adp_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyrx_adp_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyrx_adp_3 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_phyrx_adp_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module phyrx_db ( clk, srstz, x_cc, ptx_txact, r_rxdb_opt, gohi, golo, gotrans
 );
  input [1:0] r_rxdb_opt;
  input clk, srstz, x_cc, ptx_txact;
  output gohi, golo, gotrans;
  wire   N11, N12, N13, N14, N15, N16, N17, N18, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49;
  wire   [7:0] cc_buf;

  DFFQX2 cc_buf_reg_1_ ( .D(N12), .C(clk), .Q(cc_buf[1]) );
  DFFQX1 cc_buf_reg_4_ ( .D(N15), .C(clk), .Q(cc_buf[4]) );
  DFFQX1 cc_buf_reg_5_ ( .D(N16), .C(clk), .Q(cc_buf[5]) );
  DFFQX1 cc_buf_reg_6_ ( .D(N17), .C(clk), .Q(cc_buf[6]) );
  DFFQXX2 cc_buf_reg_2_ ( .D(N13), .C(clk), .Q(n4), .XQ(n3) );
  DFFQX1 cc_buf_reg_7_ ( .D(N18), .C(clk), .Q(cc_buf[7]) );
  DFFQX1 cc_buf_reg_0_ ( .D(N11), .C(clk), .Q(cc_buf[0]) );
  DFFQX1 cc_buf_reg_3_ ( .D(N14), .C(clk), .Q(cc_buf[3]) );
  XOR2X1 U3 ( .A(n26), .B(cc_buf[6]), .Y(n37) );
  NAND2X1 U4 ( .A(n6), .B(cc_buf[0]), .Y(n8) );
  NOR21XL U5 ( .B(n15), .A(n37), .Y(n14) );
  INVX2 U6 ( .A(cc_buf[1]), .Y(n25) );
  OA22X1 U7 ( .A(n31), .B(n30), .C(n29), .D(n28), .Y(n1) );
  AOI21X1 U8 ( .B(n22), .C(n21), .A(n18), .Y(n2) );
  NAND2X1 U9 ( .A(n7), .B(n8), .Y(n22) );
  NOR2X1 U10 ( .A(n22), .B(n21), .Y(n18) );
  INVX1 U11 ( .A(n3), .Y(n5) );
  NAND21X1 U12 ( .B(n1), .A(n13), .Y(n33) );
  INVX2 U13 ( .A(n24), .Y(n6) );
  NAND2X1 U14 ( .A(n24), .B(n23), .Y(n7) );
  NAND2X2 U15 ( .A(n11), .B(n10), .Y(n24) );
  AOI21X1 U16 ( .B(n14), .C(n34), .A(n32), .Y(n12) );
  INVX1 U17 ( .A(cc_buf[6]), .Y(n17) );
  INVX3 U18 ( .A(n4), .Y(n9) );
  NAND2X1 U19 ( .A(n25), .B(n9), .Y(n10) );
  NAND2X1 U20 ( .A(cc_buf[1]), .B(n4), .Y(n11) );
  XNOR2X1 U21 ( .A(n16), .B(n27), .Y(n13) );
  XOR2XL U22 ( .A(n37), .B(n36), .Y(n38) );
  INVX1 U23 ( .A(n36), .Y(n15) );
  INVXL U24 ( .A(cc_buf[7]), .Y(n21) );
  INVXL U25 ( .A(cc_buf[5]), .Y(n30) );
  INVXL U26 ( .A(cc_buf[3]), .Y(n28) );
  INVXL U27 ( .A(n20), .Y(gotrans) );
  INVX1 U28 ( .A(n44), .Y(n45) );
  INVX1 U29 ( .A(srstz), .Y(n19) );
  NAND2X1 U30 ( .A(n47), .B(n12), .Y(n44) );
  NOR21XL U31 ( .B(x_cc), .A(n19), .Y(N11) );
  INVXL U32 ( .A(cc_buf[0]), .Y(n23) );
  INVX1 U33 ( .A(n42), .Y(n43) );
  XOR2X1 U34 ( .A(n29), .B(cc_buf[3]), .Y(n36) );
  XOR2X1 U35 ( .A(n31), .B(cc_buf[5]), .Y(n29) );
  AOI21BX1 U36 ( .C(n17), .B(n2), .A(n18), .Y(n16) );
  INVX1 U37 ( .A(cc_buf[4]), .Y(n31) );
  XOR2XL U38 ( .A(n25), .B(cc_buf[0]), .Y(n20) );
  NAND21XL U39 ( .B(n25), .A(cc_buf[0]), .Y(n42) );
  NOR21XL U40 ( .B(cc_buf[3]), .A(n19), .Y(N15) );
  NOR21XL U41 ( .B(cc_buf[5]), .A(n19), .Y(N17) );
  NOR21XL U42 ( .B(cc_buf[4]), .A(n19), .Y(N16) );
  NOR21XL U43 ( .B(cc_buf[6]), .A(n19), .Y(N18) );
  AND2XL U44 ( .A(cc_buf[0]), .B(srstz), .Y(N12) );
  OAI22XL U45 ( .A(n3), .B(n25), .C(n24), .D(n23), .Y(n27) );
  NAND42X1 U46 ( .C(n5), .D(cc_buf[3]), .A(n20), .B(n42), .Y(n41) );
  AND3XL U47 ( .A(n5), .B(cc_buf[3]), .C(n43), .Y(n49) );
  AND2XL U48 ( .A(n5), .B(srstz), .Y(N14) );
  INVXL U49 ( .A(n33), .Y(n32) );
  NAND2XL U50 ( .A(n34), .B(n33), .Y(n35) );
  NAND21X2 U51 ( .B(n46), .A(n38), .Y(n39) );
  XOR2X1 U52 ( .A(n35), .B(n14), .Y(n46) );
  NAND21X2 U53 ( .B(n44), .A(n39), .Y(n40) );
  OAI22X1 U54 ( .A(n12), .B(n47), .C(n46), .D(n45), .Y(n48) );
  AO21X1 U55 ( .B(n22), .C(n21), .A(n18), .Y(n26) );
  MUX2X2 U56 ( .D0(n49), .D1(n48), .S(r_rxdb_opt[0]), .Y(gohi) );
  NAND21XL U57 ( .B(n16), .A(n27), .Y(n47) );
  NAND21X1 U58 ( .B(n13), .A(n1), .Y(n34) );
  NOR32XL U59 ( .B(cc_buf[1]), .C(srstz), .A(ptx_txact), .Y(N13) );
  MUX2IX4 U60 ( .D0(n41), .D1(n40), .S(r_rxdb_opt[1]), .Y(golo) );
endmodule


module i2cslv_a0 ( i_sda, i_scl, o_sda, i_deva, i_inc, i_fwnak, i_fwack, o_we, 
        o_re, o_r_early, o_idle, o_dec, o_busev, o_ofs, o_lt_ofs, o_wdat, 
        o_lt_buf, o_dbgpo, i_rdat, i_rd_mem, i_clk, i_rstz, i_prefetch );
  input [7:1] i_deva;
  output [3:0] o_busev;
  output [7:0] o_ofs;
  output [7:0] o_lt_ofs;
  output [7:0] o_wdat;
  output [7:0] o_lt_buf;
  output [7:0] o_dbgpo;
  input [7:0] i_rdat;
  input i_sda, i_scl, i_inc, i_fwnak, i_fwack, i_rd_mem, i_clk, i_rstz,
         i_prefetch;
  output o_sda, o_we, o_re, o_r_early, o_idle, o_dec;
  wire   i2c_scl, sdafall, cs_rwb, N74, N75, N76, N77, N78, N94, N95, N96, N97,
         N98, N99, N100, N101, N106, N107, N108, N109, N110, N111, N112, N113,
         N114, ps_rwbuf_0_, N136, N137, N138, N139, N140, N141, N142, N143,
         N144, N179, N180, N181, N182, N183, N184, N185, N186, N187, net10720,
         net10726, net10731, net10736, net10741, n61, n68, n73, n81, n97, n98,
         n99, n101, n118, n119, n120, n121, n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n62, n63, n64, n65, n66, n67,
         n69, n70, n71, n72, n74, n75, n76, n77, n78, n79, n80, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n100,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n122, n123, n124, n125, n126, n127,
         n128, n129, n130;
  wire   [1:0] cs_sta;
  wire   [7:1] add_102_carry;

  i2cdbnc_a0_1 db_scl ( .i_clk(i_clk), .i_rstz(n11), .i_i2c(i_scl), .r_opt({
        1'b1, 1'b0}), .o_i2c(i2c_scl), .rise(o_dbgpo[6]), .fall(o_dbgpo[7]) );
  i2cdbnc_a0_0 db_sda ( .i_clk(i_clk), .i_rstz(n11), .i_i2c(i_sda), .r_opt({
        1'b0, 1'b0}), .o_i2c(ps_rwbuf_0_), .rise(o_dbgpo[5]), .fall(sdafall)
         );
  SNPS_CLOCK_GATE_HIGH_i2cslv_a0_0 clk_gate_cs_bit_reg ( .CLK(i_clk), .EN(N74), 
        .ENCLK(net10720), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_i2cslv_a0_4 clk_gate_adcnt_reg ( .CLK(i_clk), .EN(N114), 
        .ENCLK(net10726), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_i2cslv_a0_3 clk_gate_rwbuf_reg ( .CLK(i_clk), .EN(N144), 
        .ENCLK(net10731), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_i2cslv_a0_2 clk_gate_lt_buf_reg ( .CLK(i_clk), .EN(N179), .ENCLK(net10736), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_i2cslv_a0_1 clk_gate_lt_ofs_reg ( .CLK(i_clk), .EN(
        o_busev[0]), .ENCLK(net10741), .TE(1'b0) );
  DFFSQX1 sdat_reg ( .D(n118), .C(i_clk), .XS(n12), .Q(o_sda) );
  DFFQX1 lt_ofs_reg_7_ ( .D(o_wdat[7]), .C(net10741), .Q(o_lt_ofs[7]) );
  DFFQX1 lt_ofs_reg_6_ ( .D(o_wdat[6]), .C(net10741), .Q(o_lt_ofs[6]) );
  DFFQX1 lt_ofs_reg_0_ ( .D(o_wdat[0]), .C(net10741), .Q(o_lt_ofs[0]) );
  DFFQX1 lt_ofs_reg_5_ ( .D(o_wdat[5]), .C(net10741), .Q(o_lt_ofs[5]) );
  DFFQX1 lt_ofs_reg_4_ ( .D(o_wdat[4]), .C(net10741), .Q(o_lt_ofs[4]) );
  DFFQX1 lt_ofs_reg_3_ ( .D(o_wdat[3]), .C(net10741), .Q(o_lt_ofs[3]) );
  DFFQX1 lt_ofs_reg_2_ ( .D(o_wdat[2]), .C(net10741), .Q(o_lt_ofs[2]) );
  DFFQX1 lt_ofs_reg_1_ ( .D(o_wdat[1]), .C(net10741), .Q(o_lt_ofs[1]) );
  DFFQX1 lt_buf_reg_7_ ( .D(N187), .C(net10736), .Q(o_lt_buf[7]) );
  DFFQX1 lt_buf_reg_6_ ( .D(N186), .C(net10736), .Q(o_lt_buf[6]) );
  DFFQX1 lt_buf_reg_5_ ( .D(N185), .C(net10736), .Q(o_lt_buf[5]) );
  DFFQX1 lt_buf_reg_4_ ( .D(N184), .C(net10736), .Q(o_lt_buf[4]) );
  DFFQX1 lt_buf_reg_3_ ( .D(N183), .C(net10736), .Q(o_lt_buf[3]) );
  DFFQX1 lt_buf_reg_2_ ( .D(N182), .C(net10736), .Q(o_lt_buf[2]) );
  DFFQX1 lt_buf_reg_1_ ( .D(N181), .C(net10736), .Q(o_lt_buf[1]) );
  DFFQX1 lt_buf_reg_0_ ( .D(N180), .C(net10736), .Q(o_lt_buf[0]) );
  DFFRQX1 adcnt_reg_2_ ( .D(N108), .C(net10726), .XR(n13), .Q(o_ofs[2]) );
  DFFRQX1 adcnt_reg_1_ ( .D(N107), .C(net10726), .XR(n13), .Q(o_ofs[1]) );
  DFFRQX1 adcnt_reg_3_ ( .D(N109), .C(net10726), .XR(n13), .Q(o_ofs[3]) );
  DFFRQX1 adcnt_reg_4_ ( .D(N110), .C(net10726), .XR(n13), .Q(o_ofs[4]) );
  DFFRQX1 adcnt_reg_5_ ( .D(N111), .C(net10726), .XR(n13), .Q(o_ofs[5]) );
  DFFRQX1 adcnt_reg_6_ ( .D(N112), .C(net10726), .XR(n14), .Q(o_ofs[6]) );
  DFFRQX1 adcnt_reg_0_ ( .D(N106), .C(net10726), .XR(n13), .Q(o_ofs[0]) );
  DFFRQX1 cs_rwb_reg ( .D(n119), .C(i_clk), .XR(n13), .Q(cs_rwb) );
  DFFSQX1 rwbuf_reg_0_ ( .D(N136), .C(net10731), .XS(n11), .Q(o_wdat[0]) );
  DFFSQX1 cs_bit_reg_1_ ( .D(N76), .C(net10720), .XS(n12), .Q(o_dbgpo[1]) );
  DFFSQX1 rwbuf_reg_7_ ( .D(N143), .C(net10731), .XS(n11), .Q(o_wdat[7]) );
  DFFSQX1 rwbuf_reg_5_ ( .D(N141), .C(net10731), .XS(n12), .Q(o_wdat[5]) );
  DFFSQX1 rwbuf_reg_6_ ( .D(N142), .C(net10731), .XS(n12), .Q(o_wdat[6]) );
  DFFSQX1 rwbuf_reg_1_ ( .D(N137), .C(net10731), .XS(n13), .Q(o_wdat[1]) );
  DFFSQX1 rwbuf_reg_2_ ( .D(N138), .C(net10731), .XS(n12), .Q(o_wdat[2]) );
  DFFSQX1 rwbuf_reg_3_ ( .D(N139), .C(net10731), .XS(n12), .Q(o_wdat[3]) );
  DFFSQX1 rwbuf_reg_4_ ( .D(N140), .C(net10731), .XS(n12), .Q(o_wdat[4]) );
  DFFSQX1 cs_bit_reg_0_ ( .D(N75), .C(net10720), .XS(n12), .Q(o_dbgpo[0]) );
  DFFRQX1 cs_sta_reg_1_ ( .D(n121), .C(i_clk), .XR(n14), .Q(cs_sta[1]) );
  DFFRQX1 adcnt_reg_7_ ( .D(N113), .C(net10726), .XR(n13), .Q(o_ofs[7]) );
  DFFRQX1 cs_sta_reg_0_ ( .D(n120), .C(i_clk), .XR(n13), .Q(cs_sta[0]) );
  DFFSQX1 cs_bit_reg_2_ ( .D(N77), .C(net10720), .XS(n12), .Q(o_dbgpo[2]) );
  DFFSQX1 cs_bit_reg_3_ ( .D(N78), .C(net10720), .XS(n12), .Q(o_dbgpo[3]) );
  AOI21X1 U3 ( .B(n108), .C(o_dbgpo[7]), .A(n90), .Y(n1) );
  INVX1 U4 ( .A(n57), .Y(n2) );
  GEN2XL U5 ( .D(n116), .E(n30), .C(n108), .B(o_dbgpo[7]), .A(o_busev[0]), .Y(
        N114) );
  INVX1 U6 ( .A(n15), .Y(n12) );
  INVX1 U7 ( .A(n15), .Y(n13) );
  INVX1 U8 ( .A(n15), .Y(n14) );
  XNOR2XL U9 ( .A(i_fwnak), .B(i_fwack), .Y(n61) );
  INVX1 U10 ( .A(n15), .Y(n11) );
  INVX1 U11 ( .A(i_rstz), .Y(n15) );
  INVX1 U12 ( .A(n69), .Y(n93) );
  INVX1 U13 ( .A(o_dbgpo[7]), .Y(n125) );
  INVX1 U14 ( .A(n112), .Y(n49) );
  INVX1 U15 ( .A(n81), .Y(n100) );
  INVX1 U16 ( .A(n98), .Y(n122) );
  AND2X1 U17 ( .A(n2), .B(n106), .Y(o_dec) );
  NAND21X1 U18 ( .B(n85), .A(o_busev[1]), .Y(n34) );
  INVX1 U19 ( .A(n25), .Y(o_busev[1]) );
  NAND32X1 U20 ( .B(n54), .C(n26), .A(n108), .Y(n25) );
  INVX1 U21 ( .A(o_dbgpo[6]), .Y(n26) );
  NAND21X1 U22 ( .B(n54), .A(i_prefetch), .Y(n112) );
  INVX1 U23 ( .A(n57), .Y(n108) );
  AND4X1 U24 ( .A(n109), .B(o_dbgpo[6]), .C(n108), .D(n107), .Y(n111) );
  INVX1 U25 ( .A(n18), .Y(n17) );
  INVX1 U26 ( .A(n83), .Y(n107) );
  INVX1 U27 ( .A(n114), .Y(n109) );
  INVX1 U28 ( .A(n35), .Y(o_we) );
  INVX1 U29 ( .A(n27), .Y(n116) );
  GEN2XL U30 ( .D(n124), .E(i_fwnak), .C(n64), .B(n125), .A(n63), .Y(n118) );
  INVX1 U31 ( .A(n61), .Y(n124) );
  AND3X1 U32 ( .A(n61), .B(i_rdat[7]), .C(n36), .Y(n64) );
  MUX2X1 U33 ( .D0(n62), .D1(n60), .S(n125), .Y(n63) );
  INVX1 U34 ( .A(i_rd_mem), .Y(n123) );
  NAND32X1 U35 ( .B(n26), .C(n92), .A(n76), .Y(n69) );
  AO22AXL U36 ( .A(i_rdat[3]), .B(n92), .C(n93), .D(n130), .Y(N139) );
  AO22AXL U37 ( .A(i_rdat[2]), .B(n92), .C(n93), .D(n127), .Y(N138) );
  AO22X1 U38 ( .A(n93), .B(o_wdat[0]), .C(i_rdat[1]), .D(n92), .Y(N137) );
  OA21X1 U39 ( .B(n93), .C(n92), .A(n70), .Y(N144) );
  ENOX1 U40 ( .A(n69), .B(n67), .C(n92), .D(i_rdat[7]), .Y(N143) );
  INVX1 U41 ( .A(n59), .Y(n36) );
  INVX1 U42 ( .A(n19), .Y(o_busev[0]) );
  NAND32X1 U43 ( .B(n125), .C(n65), .A(n51), .Y(n19) );
  INVX1 U44 ( .A(n54), .Y(n51) );
  INVX1 U45 ( .A(n73), .Y(o_busev[2]) );
  OR2X1 U46 ( .A(n100), .B(n3), .Y(n96) );
  AOI21X1 U47 ( .B(n86), .C(n85), .A(n88), .Y(n3) );
  GEN2XL U48 ( .D(n89), .E(o_dbgpo[7]), .C(n88), .B(n106), .A(n100), .Y(n90)
         );
  INVX1 U49 ( .A(i_prefetch), .Y(n82) );
  INVX1 U50 ( .A(n76), .Y(n106) );
  NOR2X1 U51 ( .A(o_busev[3]), .B(o_busev[2]), .Y(n81) );
  INVX1 U52 ( .A(n84), .Y(n88) );
  NAND5XL U53 ( .A(n125), .B(o_dbgpo[6]), .C(n108), .D(n83), .E(n82), .Y(n84)
         );
  NAND32X1 U54 ( .B(n72), .C(n125), .A(n71), .Y(n97) );
  INVX1 U55 ( .A(o_idle), .Y(n71) );
  INVX1 U56 ( .A(n70), .Y(n72) );
  INVX1 U57 ( .A(n77), .Y(n80) );
  NAND21X1 U58 ( .B(n97), .A(n76), .Y(n77) );
  GEN2XL U59 ( .D(n75), .E(o_dbgpo[3]), .C(n106), .B(n74), .A(n78), .Y(N78) );
  INVX1 U60 ( .A(n99), .Y(n75) );
  INVX1 U61 ( .A(n97), .Y(n74) );
  NAND2X1 U62 ( .A(n34), .B(n35), .Y(N179) );
  NAND2X1 U63 ( .A(n73), .B(n98), .Y(n78) );
  AO21X1 U64 ( .B(o_we), .C(o_wdat[0]), .A(n110), .Y(N180) );
  AO21X1 U65 ( .B(n80), .C(n79), .A(n78), .Y(N75) );
  NAND2X1 U66 ( .A(o_busev[3]), .B(n73), .Y(n98) );
  OAI22X1 U67 ( .A(n33), .B(n35), .C(n34), .D(n32), .Y(N184) );
  OAI22X1 U68 ( .A(n39), .B(n35), .C(n34), .D(n33), .Y(N185) );
  OAI22X1 U69 ( .A(n67), .B(n35), .C(n34), .D(n39), .Y(N186) );
  OAI22X1 U70 ( .A(n127), .B(n35), .C(n126), .D(n34), .Y(N181) );
  OAI22X1 U71 ( .A(n130), .B(n35), .C(n127), .D(n34), .Y(N182) );
  OAI22X1 U72 ( .A(n32), .B(n35), .C(n130), .D(n34), .Y(N183) );
  NAND3X1 U73 ( .A(n97), .B(n73), .C(n98), .Y(N74) );
  INVX1 U74 ( .A(n101), .Y(n128) );
  INVX1 U75 ( .A(n65), .Y(n66) );
  BUFX3 U76 ( .A(o_busev[3]), .Y(o_dbgpo[4]) );
  NOR43XL U77 ( .B(n23), .C(n22), .D(n21), .A(n20), .Y(n24) );
  XOR2X1 U78 ( .A(i_deva[5]), .B(o_wdat[4]), .Y(n20) );
  XOR2X1 U79 ( .A(n37), .B(o_wdat[5]), .Y(n23) );
  XOR2X1 U80 ( .A(n40), .B(o_wdat[6]), .Y(n21) );
  NAND21X1 U81 ( .B(n18), .A(o_dbgpo[0]), .Y(n54) );
  OR3XL U82 ( .A(o_dbgpo[2]), .B(o_dbgpo[3]), .C(o_dbgpo[1]), .Y(n18) );
  NAND4X1 U83 ( .A(n4), .B(n5), .C(n6), .D(n24), .Y(n85) );
  XNOR2XL U84 ( .A(o_wdat[1]), .B(i_deva[2]), .Y(n4) );
  XNOR2XL U85 ( .A(o_wdat[0]), .B(i_deva[1]), .Y(n5) );
  XNOR2XL U86 ( .A(o_wdat[2]), .B(i_deva[3]), .Y(n6) );
  XOR2X1 U87 ( .A(n38), .B(o_wdat[3]), .Y(n22) );
  AND3X1 U88 ( .A(o_dbgpo[6]), .B(n116), .C(n115), .Y(o_re) );
  MUX2X1 U89 ( .D0(n111), .D1(n110), .S(i_prefetch), .Y(o_r_early) );
  OAI32X1 U90 ( .A(i_prefetch), .B(ps_rwbuf_0_), .C(n114), .D(n113), .E(n112), 
        .Y(n115) );
  INVX1 U91 ( .A(n31), .Y(n110) );
  NAND21X1 U92 ( .B(n34), .A(ps_rwbuf_0_), .Y(n31) );
  INVX1 U93 ( .A(i_deva[4]), .Y(n38) );
  NAND21X1 U94 ( .B(o_dbgpo[0]), .A(n17), .Y(n76) );
  NAND43X1 U95 ( .B(n48), .C(n47), .D(n46), .A(n45), .Y(n83) );
  XOR2X1 U96 ( .A(o_wdat[2]), .B(i_deva[2]), .Y(n48) );
  XOR2X1 U97 ( .A(i_deva[1]), .B(o_wdat[1]), .Y(n47) );
  AND4X1 U98 ( .A(n44), .B(n43), .C(n42), .D(n41), .Y(n45) );
  NAND21X1 U99 ( .B(n76), .A(cs_rwb), .Y(n114) );
  NAND21X1 U100 ( .B(cs_sta[0]), .A(n89), .Y(n57) );
  XOR2X1 U101 ( .A(n40), .B(o_wdat[7]), .Y(n41) );
  XOR2X1 U102 ( .A(n39), .B(i_deva[5]), .Y(n42) );
  XOR2X1 U103 ( .A(n37), .B(o_wdat[6]), .Y(n44) );
  XOR2X1 U104 ( .A(n38), .B(o_wdat[4]), .Y(n43) );
  XOR2X1 U105 ( .A(i_deva[3]), .B(o_wdat[3]), .Y(n46) );
  INVX1 U106 ( .A(cs_sta[1]), .Y(n89) );
  INVX1 U107 ( .A(o_wdat[5]), .Y(n39) );
  INVX1 U108 ( .A(i_deva[7]), .Y(n40) );
  INVX1 U109 ( .A(i_deva[6]), .Y(n37) );
  NAND43X1 U110 ( .B(cs_rwb), .C(n27), .D(n54), .A(o_dbgpo[7]), .Y(n35) );
  NAND21X1 U111 ( .B(cs_sta[0]), .A(cs_sta[1]), .Y(n27) );
  INVX1 U112 ( .A(cs_rwb), .Y(n113) );
  AOI22X1 U113 ( .A(i_rd_mem), .B(i_rdat[7]), .C(n123), .D(o_wdat[7]), .Y(n68)
         );
  AO21X1 U114 ( .B(ps_rwbuf_0_), .C(n106), .A(n53), .Y(n55) );
  MUX2X1 U115 ( .D0(n52), .D1(cs_rwb), .S(n51), .Y(n53) );
  NAND21X1 U116 ( .B(n117), .A(cs_rwb), .Y(n52) );
  INVX1 U117 ( .A(n68), .Y(n117) );
  OAI211X1 U118 ( .C(n58), .D(n57), .A(n70), .B(n56), .Y(n62) );
  MUX2X1 U119 ( .D0(n50), .D1(n68), .S(n109), .Y(n58) );
  AOI22X1 U120 ( .A(cs_sta[1]), .B(n55), .C(cs_sta[0]), .D(n54), .Y(n56) );
  AO21X1 U121 ( .B(n107), .C(n51), .A(n49), .Y(n50) );
  AND4X1 U122 ( .A(o_dbgpo[2]), .B(o_dbgpo[1]), .C(o_dbgpo[3]), .D(o_dbgpo[0]), 
        .Y(o_idle) );
  NAND2X1 U123 ( .A(n7), .B(n59), .Y(n92) );
  NAND4X1 U124 ( .A(cs_rwb), .B(n17), .C(n70), .D(i_rd_mem), .Y(n7) );
  NAND6XL U125 ( .A(n99), .B(cs_rwb), .C(n70), .D(n16), .E(i_rd_mem), .F(
        o_dbgpo[3]), .Y(n59) );
  INVX1 U126 ( .A(i2c_scl), .Y(n16) );
  AO22X1 U127 ( .A(o_wdat[5]), .B(n93), .C(i_rdat[6]), .D(n92), .Y(N142) );
  AO22X1 U128 ( .A(o_wdat[4]), .B(n93), .C(i_rdat[5]), .D(n92), .Y(N141) );
  AO22X1 U129 ( .A(o_wdat[3]), .B(n93), .C(i_rdat[4]), .D(n92), .Y(N140) );
  AND3X1 U130 ( .A(o_sda), .B(n61), .C(n59), .Y(n60) );
  OAI21BBX1 U131 ( .A(i_rdat[0]), .B(n92), .C(n8), .Y(N136) );
  NAND4X1 U132 ( .A(ps_rwbuf_0_), .B(o_dbgpo[6]), .C(n76), .D(n113), .Y(n8) );
  NOR32XL U133 ( .B(i2c_scl), .C(o_dbgpo[5]), .A(o_dbgpo[7]), .Y(o_busev[3])
         );
  NAND3X1 U134 ( .A(i2c_scl), .B(n125), .C(sdafall), .Y(n73) );
  AO222X1 U135 ( .A(o_ofs[6]), .B(n108), .C(N100), .D(n116), .E(o_wdat[6]), 
        .F(n66), .Y(N112) );
  NAND21X1 U136 ( .B(cs_sta[1]), .A(cs_sta[0]), .Y(n65) );
  AO222X1 U137 ( .A(o_ofs[7]), .B(n108), .C(N101), .D(n116), .E(o_wdat[7]), 
        .F(n66), .Y(N113) );
  MUX2X1 U138 ( .D0(n91), .D1(cs_sta[0]), .S(n1), .Y(n120) );
  NAND21X1 U139 ( .B(n87), .A(n96), .Y(n91) );
  AND4X1 U140 ( .A(n81), .B(n106), .C(n113), .D(n102), .Y(n87) );
  MUX2X1 U141 ( .D0(n105), .D1(cs_sta[1]), .S(n1), .Y(n121) );
  NAND21X1 U142 ( .B(n104), .A(n103), .Y(n105) );
  AO21X1 U143 ( .B(n114), .C(n102), .A(n100), .Y(n103) );
  INVX1 U144 ( .A(n96), .Y(n104) );
  AO222X1 U145 ( .A(o_ofs[5]), .B(n108), .C(N99), .D(n116), .E(o_wdat[5]), .F(
        n66), .Y(N111) );
  AO222X1 U146 ( .A(o_ofs[4]), .B(n108), .C(N98), .D(n116), .E(o_wdat[4]), .F(
        n66), .Y(N110) );
  AO222X1 U147 ( .A(o_ofs[3]), .B(n108), .C(N97), .D(n116), .E(o_wdat[3]), .F(
        n66), .Y(N109) );
  NAND21X1 U148 ( .B(n89), .A(cs_sta[0]), .Y(n70) );
  GEN2XL U149 ( .D(n128), .E(o_dbgpo[2]), .C(n99), .B(n80), .A(n122), .Y(N77)
         );
  GEN2XL U150 ( .D(o_dbgpo[1]), .E(o_dbgpo[0]), .C(n101), .B(n80), .A(n122), 
        .Y(N76) );
  MUX2BXL U151 ( .D0(n106), .D1(n9), .S(cs_rwb), .Y(n30) );
  AOI21X1 U152 ( .B(n51), .C(n82), .A(n86), .Y(n9) );
  MUX2X1 U153 ( .D0(n95), .D1(ps_rwbuf_0_), .S(n94), .Y(n119) );
  AND2X1 U154 ( .A(n73), .B(o_busev[1]), .Y(n94) );
  AND2X1 U155 ( .A(cs_rwb), .B(n73), .Y(n95) );
  NOR2X1 U156 ( .A(n128), .B(o_dbgpo[2]), .Y(n99) );
  NOR2X1 U157 ( .A(o_dbgpo[1]), .B(o_dbgpo[0]), .Y(n101) );
  OAI22AX1 U158 ( .D(o_wdat[7]), .C(n35), .A(n34), .B(n67), .Y(N187) );
  INVX1 U159 ( .A(n29), .Y(n86) );
  NAND5XL U160 ( .A(o_dbgpo[1]), .B(i_prefetch), .C(n129), .D(n28), .E(n79), 
        .Y(n29) );
  INVX1 U161 ( .A(o_dbgpo[2]), .Y(n28) );
  INVX1 U162 ( .A(o_dbgpo[0]), .Y(n79) );
  INVX1 U163 ( .A(o_dbgpo[3]), .Y(n129) );
  AO222X1 U164 ( .A(o_ofs[2]), .B(n2), .C(N96), .D(n116), .E(o_wdat[2]), .F(
        n66), .Y(N108) );
  AO222X1 U165 ( .A(o_ofs[1]), .B(n2), .C(N95), .D(n116), .E(o_wdat[1]), .F(
        n66), .Y(N107) );
  AO222X1 U166 ( .A(o_ofs[0]), .B(n2), .C(N94), .D(n116), .E(o_wdat[0]), .F(
        n66), .Y(N106) );
  INVX1 U167 ( .A(cs_sta[0]), .Y(n102) );
  INVX1 U168 ( .A(o_wdat[2]), .Y(n130) );
  INVX1 U169 ( .A(o_wdat[1]), .Y(n127) );
  INVX1 U170 ( .A(o_wdat[0]), .Y(n126) );
  INVX1 U171 ( .A(o_wdat[6]), .Y(n67) );
  INVX1 U172 ( .A(o_wdat[3]), .Y(n32) );
  INVX1 U173 ( .A(o_wdat[4]), .Y(n33) );
  XOR2X1 U174 ( .A(o_ofs[7]), .B(add_102_carry[7]), .Y(N101) );
  AND2X1 U175 ( .A(o_ofs[6]), .B(add_102_carry[6]), .Y(add_102_carry[7]) );
  XOR2X1 U176 ( .A(add_102_carry[6]), .B(o_ofs[6]), .Y(N100) );
  AND2X1 U177 ( .A(o_ofs[5]), .B(add_102_carry[5]), .Y(add_102_carry[6]) );
  XOR2X1 U178 ( .A(add_102_carry[5]), .B(o_ofs[5]), .Y(N99) );
  AND2X1 U179 ( .A(o_ofs[4]), .B(add_102_carry[4]), .Y(add_102_carry[5]) );
  XOR2X1 U180 ( .A(add_102_carry[4]), .B(o_ofs[4]), .Y(N98) );
  AND2X1 U181 ( .A(o_ofs[3]), .B(add_102_carry[3]), .Y(add_102_carry[4]) );
  XOR2X1 U182 ( .A(add_102_carry[3]), .B(o_ofs[3]), .Y(N97) );
  AND2X1 U183 ( .A(o_ofs[2]), .B(add_102_carry[2]), .Y(add_102_carry[3]) );
  XOR2X1 U184 ( .A(add_102_carry[2]), .B(o_ofs[2]), .Y(N96) );
  AND2X1 U185 ( .A(o_ofs[1]), .B(add_102_carry[1]), .Y(add_102_carry[2]) );
  XOR2X1 U186 ( .A(add_102_carry[1]), .B(o_ofs[1]), .Y(N95) );
  AND2X1 U187 ( .A(i_inc), .B(o_ofs[0]), .Y(add_102_carry[1]) );
  XOR2X1 U188 ( .A(o_ofs[0]), .B(i_inc), .Y(N94) );
endmodule


module SNPS_CLOCK_GATE_HIGH_i2cslv_a0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_i2cslv_a0_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_i2cslv_a0_3 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_i2cslv_a0_4 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_i2cslv_a0_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module i2cdbnc_a0_0 ( i_clk, i_rstz, i_i2c, r_opt, o_i2c, rise, fall );
  input [1:0] r_opt;
  input i_clk, i_rstz, i_i2c;
  output o_i2c, rise, fall;
  wire   d_i2c_2_, N18, N19, n2, n7, n8, n9, n10, n11;

  DFFSQX1 d_i2c_reg_2_ ( .D(N19), .C(i_clk), .XS(i_rstz), .Q(d_i2c_2_) );
  DFFSQX1 d_i2c_reg_0_ ( .D(i_i2c), .C(i_clk), .XS(i_rstz), .Q(N18) );
  DFFSQX1 d_i2c_reg_1_ ( .D(N18), .C(i_clk), .XS(i_rstz), .Q(N19) );
  DFFSQXX1 r_i2c_reg ( .D(n7), .C(i_clk), .XS(i_rstz), .Q(o_i2c), .XQ(n11) );
  INVX1 U3 ( .A(n10), .Y(rise) );
  OAI211X1 U4 ( .C(d_i2c_2_), .D(r_opt[0]), .A(n11), .B(n9), .Y(n10) );
  AND2X1 U5 ( .A(N18), .B(N19), .Y(n9) );
  AOI211X1 U6 ( .C(n2), .D(d_i2c_2_), .A(n11), .B(n8), .Y(fall) );
  INVX1 U7 ( .A(r_opt[1]), .Y(n2) );
  OR2X1 U8 ( .A(N19), .B(N18), .Y(n8) );
  OAI21X1 U9 ( .B(fall), .C(n11), .A(n10), .Y(n7) );
endmodule


module i2cdbnc_a0_1 ( i_clk, i_rstz, i_i2c, r_opt, o_i2c, rise, fall );
  input [1:0] r_opt;
  input i_clk, i_rstz, i_i2c;
  output o_i2c, rise, fall;
  wire   d_i2c_2_, N18, N19, n1, n6, n2, n3, n4, n5;

  DFFSQX1 d_i2c_reg_0_ ( .D(i_i2c), .C(i_clk), .XS(i_rstz), .Q(N18) );
  DFFSQX1 d_i2c_reg_1_ ( .D(N18), .C(i_clk), .XS(i_rstz), .Q(N19) );
  DFFSQX1 d_i2c_reg_2_ ( .D(N19), .C(i_clk), .XS(i_rstz), .Q(d_i2c_2_) );
  DFFSQXXL r_i2c_reg ( .D(n6), .C(i_clk), .XS(i_rstz), .Q(o_i2c), .XQ(n1) );
  INVX1 U3 ( .A(n5), .Y(fall) );
  AO21X1 U4 ( .B(n5), .C(o_i2c), .A(rise), .Y(n6) );
  NOR43XL U5 ( .B(n1), .C(N19), .D(N18), .A(n4), .Y(rise) );
  NOR2X1 U6 ( .A(d_i2c_2_), .B(r_opt[0]), .Y(n4) );
  NAND32X1 U7 ( .B(N19), .C(N18), .A(n3), .Y(n5) );
  OA21X1 U8 ( .B(r_opt[1]), .C(n2), .A(o_i2c), .Y(n3) );
  INVX1 U9 ( .A(d_i2c_2_), .Y(n2) );
endmodule


module regbank_a0 ( srci, dm_fault, cc1_di, cc2_di, di_rd_det, di_stbovp, 
        i_tmrf, i_vcbyval, dnchk_en, r_pwrv_upd, aswkup, ps_pwrdn, r_sleep, 
        r_pwrdn, r_ocdrv_enz, r_osc_stop, r_osc_lo, r_osc_gate, r_fw_pwrv, 
        r_cvcwr, r_cvofs, r_otpi_gate, r_pwrctl, r_pwr_i, r_cvctl, r_srcctl, 
        r_dpdmctl, r_ccrx, r_cctrx, r_ccctl, r_fcpwr, r_fcpre, fcp_r_dat, 
        fcp_r_sta, fcp_r_msk, fcp_r_ctl, fcp_r_crc, fcp_r_acc, fcp_r_tui, 
        r_accctl, r_bclk_sel, r_dacwr, r_dac_en, r_sar_en, r_adofs, r_isofs, 
        x_daclsb, r_comp_opt, dac_r_ctl, dac_r_comp, dac_r_cmpsta, dac_r_vs, 
        REVID, atpg_en, sfr_r, sfr_w, set_hold, bkpt_hold, cpurst, sfr_addr, 
        sfr_wdat, sfr_rdat, ff_p0, di_p0, ictlr_idle, ictlr_inc, r_inst_ofs, 
        r_psrd, r_pswr, r_fortxdat, r_fortxrdy, r_fortxen, r_ana_tm, r_gpio_tm, 
        r_gpio_ie, r_gpio_oe, r_gpio_pu, r_gpio_pd, r_gpio_s0, r_gpio_s1, 
        r_gpio_s2, r_gpio_s3, r_regtrm, i_pc, i_goidle, i_gobusy, i_i2c_idle, 
        bus_idle, i2c_stretch, i_i2c_rwbuf, i_i2c_ltbuf, i_i2c_ofs, o_intr, 
        r_auto_gdcrc, r_exist1st, r_ordrs4, r_fifopsh, r_fifopop, r_unlock, 
        r_first, r_last, r_fiforst, r_set_cpmsgid, r_txendk, r_txnumk, 
        r_txshrt, r_auto_discard, r_hold_mcu, r_txauto, r_rxords_ena, r_spec, 
        r_dat_spec, r_dat_portrole, r_dat_datarole, r_discard, r_pshords, 
        r_pg0_sel, r_strtch, r_i2c_attr, r_i2c_ninc, r_hwi2c_en, r_i2c_fwnak, 
        r_i2c_fwack, r_i2c_deva, i2c_ev, prl_c0set, prl_cany0, prl_discard, 
        prl_GCTxDone, prl_cpmsgid, pff_ack, prx_rst, pff_obsd, pff_full, 
        pff_empty, ptx_ack, pff_ptr, prx_adpn, pff_rdat, pff_rxpart, 
        prx_rcvinf, ptx_fsm, prx_fsm, prl_fsm, prx_setsta, clk_1500k, clk_500k, 
        clk_500, clk, xrstz, xclk, dbgpo, srstz, prstz );
  input [5:0] srci;
  output [11:0] r_fw_pwrv;
  output [1:0] r_cvcwr;
  input [15:0] r_cvofs;
  output [7:4] r_pwrctl;
  output [7:0] r_pwr_i;
  output [7:0] r_cvctl;
  output [7:0] r_srcctl;
  output [7:0] r_dpdmctl;
  output [7:0] r_ccrx;
  output [7:0] r_cctrx;
  output [7:0] r_ccctl;
  output [6:0] r_fcpwr;
  input [7:0] fcp_r_dat;
  input [7:0] fcp_r_sta;
  input [7:0] fcp_r_msk;
  input [7:0] fcp_r_ctl;
  input [7:0] fcp_r_crc;
  input [7:0] fcp_r_acc;
  input [7:0] fcp_r_tui;
  input [7:0] r_accctl;
  output [14:0] r_dacwr;
  input [7:0] r_dac_en;
  input [7:0] r_sar_en;
  input [7:0] r_adofs;
  input [7:0] r_isofs;
  input [5:0] x_daclsb;
  output [7:0] r_comp_opt;
  input [7:0] dac_r_ctl;
  input [7:0] dac_r_comp;
  input [7:0] dac_r_cmpsta;
  input [63:0] dac_r_vs;
  input [6:0] REVID;
  input [7:0] sfr_addr;
  input [7:0] sfr_wdat;
  output [7:0] sfr_rdat;
  input [7:0] ff_p0;
  input [7:0] di_p0;
  output [14:0] r_inst_ofs;
  output [3:0] r_ana_tm;
  output [1:0] r_gpio_ie;
  output [6:0] r_gpio_oe;
  output [6:0] r_gpio_pu;
  output [6:0] r_gpio_pd;
  output [2:0] r_gpio_s0;
  output [2:0] r_gpio_s1;
  output [2:0] r_gpio_s2;
  output [2:0] r_gpio_s3;
  output [55:0] r_regtrm;
  input [15:0] i_pc;
  input [7:0] i_i2c_rwbuf;
  input [7:0] i_i2c_ltbuf;
  input [7:0] i_i2c_ofs;
  output [4:0] o_intr;
  output [1:0] r_auto_gdcrc;
  output [4:0] r_txnumk;
  output [6:0] r_txauto;
  output [6:0] r_rxords_ena;
  output [1:0] r_spec;
  output [1:0] r_dat_spec;
  output [3:0] r_pg0_sel;
  output [7:1] r_i2c_deva;
  input [7:0] i2c_ev;
  input [2:0] prl_cpmsgid;
  input [1:0] pff_ack;
  input [1:0] prx_rst;
  input [5:0] pff_ptr;
  input [5:0] prx_adpn;
  input [7:0] pff_rdat;
  input [15:0] pff_rxpart;
  input [4:0] prx_rcvinf;
  input [2:0] ptx_fsm;
  input [3:0] prx_fsm;
  input [3:0] prl_fsm;
  input [6:0] prx_setsta;
  output [31:0] dbgpo;
  input dm_fault, cc1_di, cc2_di, di_rd_det, di_stbovp, i_tmrf, i_vcbyval,
         dnchk_en, atpg_en, sfr_r, sfr_w, set_hold, bkpt_hold, cpurst,
         ictlr_idle, ictlr_inc, i_goidle, i_gobusy, i_i2c_idle, prl_c0set,
         prl_cany0, prl_discard, prl_GCTxDone, pff_obsd, pff_full, pff_empty,
         ptx_ack, clk_1500k, clk_500k, clk_500, clk, xrstz, xclk;
  output r_pwrv_upd, aswkup, ps_pwrdn, r_sleep, r_pwrdn, r_ocdrv_enz,
         r_osc_stop, r_osc_lo, r_osc_gate, r_otpi_gate, r_fcpre, r_bclk_sel,
         r_psrd, r_pswr, r_fortxdat, r_fortxrdy, r_fortxen, r_gpio_tm,
         bus_idle, i2c_stretch, r_exist1st, r_ordrs4, r_fifopsh, r_fifopop,
         r_unlock, r_first, r_last, r_fiforst, r_set_cpmsgid, r_txendk,
         r_txshrt, r_auto_discard, r_hold_mcu, r_dat_portrole, r_dat_datarole,
         r_discard, r_pshords, r_strtch, r_i2c_attr, r_i2c_ninc, r_hwi2c_en,
         r_i2c_fwnak, r_i2c_fwack, srstz, prstz;
  wire   hit_223, hit_207, hit_206, hit_202, hit_201, hit_197, hit_195,
         hit_194, hit_151, we_246, we_245, we_232, we_231, we_230, we_228,
         we_227, we_222, we_217, we_215, we_214, we_213, we_211, we_209,
         we_203, we_191, we_187, we_182, we_181, we_176, we_175, we_172,
         we_171, we_148, we_143, regF4_7_, regF4_3, regE3_0, regD3_7_, regD3_3,
         reg25_0_, reg19_7_, reg12_1, reg11_7_, reg11_4, regAD_7, N23, N24,
         N25, N26, N27, N29, N30, N31, N32, N33, N34, N35, N36, upd01, phyrst,
         upd12, upd18, upd19, upd20, upd21, lt_reg26_0, i2c_mode_upd,
         i2c_mode_wdat, upd31, N81, as_p0_chg, dmf_wkup, p0_chg_clr,
         di_stbovp_clr, di_rd_det_clr, dm_fault_clr, pwrdn_rstz, osc_low_clr,
         osc_low_rstz, r_pos_gate, m_ovp, m_ovp_sta, setAE_7, m_scp, m_scp_sta,
         s_ovp, s_ovp_sta, s_scp, s_scp_sta, net10758, n1076, n1095, n1096,
         n1120, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
         n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
         n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, SYNOPSYS_UNCONNECTED_1,
         SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3,
         SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5,
         SYNOPSYS_UNCONNECTED_6, SYNOPSYS_UNCONNECTED_7,
         SYNOPSYS_UNCONNECTED_8, SYNOPSYS_UNCONNECTED_9,
         SYNOPSYS_UNCONNECTED_10, SYNOPSYS_UNCONNECTED_11,
         SYNOPSYS_UNCONNECTED_12, SYNOPSYS_UNCONNECTED_13,
         SYNOPSYS_UNCONNECTED_14, SYNOPSYS_UNCONNECTED_15,
         SYNOPSYS_UNCONNECTED_16, SYNOPSYS_UNCONNECTED_17,
         SYNOPSYS_UNCONNECTED_18, SYNOPSYS_UNCONNECTED_19,
         SYNOPSYS_UNCONNECTED_20, SYNOPSYS_UNCONNECTED_21,
         SYNOPSYS_UNCONNECTED_22, SYNOPSYS_UNCONNECTED_23,
         SYNOPSYS_UNCONNECTED_24, SYNOPSYS_UNCONNECTED_25,
         SYNOPSYS_UNCONNECTED_26, SYNOPSYS_UNCONNECTED_27,
         SYNOPSYS_UNCONNECTED_28, SYNOPSYS_UNCONNECTED_29,
         SYNOPSYS_UNCONNECTED_30, SYNOPSYS_UNCONNECTED_31,
         SYNOPSYS_UNCONNECTED_32, SYNOPSYS_UNCONNECTED_33,
         SYNOPSYS_UNCONNECTED_34, SYNOPSYS_UNCONNECTED_35,
         SYNOPSYS_UNCONNECTED_36, SYNOPSYS_UNCONNECTED_37,
         SYNOPSYS_UNCONNECTED_38, SYNOPSYS_UNCONNECTED_39,
         SYNOPSYS_UNCONNECTED_40, SYNOPSYS_UNCONNECTED_41,
         SYNOPSYS_UNCONNECTED_42, SYNOPSYS_UNCONNECTED_43,
         SYNOPSYS_UNCONNECTED_44, SYNOPSYS_UNCONNECTED_45,
         SYNOPSYS_UNCONNECTED_46, SYNOPSYS_UNCONNECTED_47,
         SYNOPSYS_UNCONNECTED_48, SYNOPSYS_UNCONNECTED_49,
         SYNOPSYS_UNCONNECTED_50, SYNOPSYS_UNCONNECTED_51,
         SYNOPSYS_UNCONNECTED_52, SYNOPSYS_UNCONNECTED_53,
         SYNOPSYS_UNCONNECTED_54, SYNOPSYS_UNCONNECTED_55,
         SYNOPSYS_UNCONNECTED_56, SYNOPSYS_UNCONNECTED_57,
         SYNOPSYS_UNCONNECTED_58, SYNOPSYS_UNCONNECTED_59,
         SYNOPSYS_UNCONNECTED_60, SYNOPSYS_UNCONNECTED_61,
         SYNOPSYS_UNCONNECTED_62, SYNOPSYS_UNCONNECTED_63,
         SYNOPSYS_UNCONNECTED_64, SYNOPSYS_UNCONNECTED_65,
         SYNOPSYS_UNCONNECTED_66, SYNOPSYS_UNCONNECTED_67,
         SYNOPSYS_UNCONNECTED_68, SYNOPSYS_UNCONNECTED_69,
         SYNOPSYS_UNCONNECTED_70, SYNOPSYS_UNCONNECTED_71,
         SYNOPSYS_UNCONNECTED_72, SYNOPSYS_UNCONNECTED_73,
         SYNOPSYS_UNCONNECTED_74, SYNOPSYS_UNCONNECTED_75,
         SYNOPSYS_UNCONNECTED_76, SYNOPSYS_UNCONNECTED_77,
         SYNOPSYS_UNCONNECTED_78, SYNOPSYS_UNCONNECTED_79,
         SYNOPSYS_UNCONNECTED_80, SYNOPSYS_UNCONNECTED_81,
         SYNOPSYS_UNCONNECTED_82, SYNOPSYS_UNCONNECTED_83,
         SYNOPSYS_UNCONNECTED_84, SYNOPSYS_UNCONNECTED_85,
         SYNOPSYS_UNCONNECTED_86, SYNOPSYS_UNCONNECTED_87,
         SYNOPSYS_UNCONNECTED_88, SYNOPSYS_UNCONNECTED_89,
         SYNOPSYS_UNCONNECTED_90, SYNOPSYS_UNCONNECTED_91,
         SYNOPSYS_UNCONNECTED_92, SYNOPSYS_UNCONNECTED_93,
         SYNOPSYS_UNCONNECTED_94, SYNOPSYS_UNCONNECTED_95,
         SYNOPSYS_UNCONNECTED_96, SYNOPSYS_UNCONNECTED_97,
         SYNOPSYS_UNCONNECTED_98, SYNOPSYS_UNCONNECTED_99,
         SYNOPSYS_UNCONNECTED_100, SYNOPSYS_UNCONNECTED_101,
         SYNOPSYS_UNCONNECTED_102, SYNOPSYS_UNCONNECTED_103,
         SYNOPSYS_UNCONNECTED_104, SYNOPSYS_UNCONNECTED_105,
         SYNOPSYS_UNCONNECTED_106, SYNOPSYS_UNCONNECTED_107,
         SYNOPSYS_UNCONNECTED_108, SYNOPSYS_UNCONNECTED_109,
         SYNOPSYS_UNCONNECTED_110, SYNOPSYS_UNCONNECTED_111,
         SYNOPSYS_UNCONNECTED_112, SYNOPSYS_UNCONNECTED_113,
         SYNOPSYS_UNCONNECTED_114, SYNOPSYS_UNCONNECTED_115,
         SYNOPSYS_UNCONNECTED_116, SYNOPSYS_UNCONNECTED_117,
         SYNOPSYS_UNCONNECTED_118, SYNOPSYS_UNCONNECTED_119,
         SYNOPSYS_UNCONNECTED_120, SYNOPSYS_UNCONNECTED_121,
         SYNOPSYS_UNCONNECTED_122, SYNOPSYS_UNCONNECTED_123,
         SYNOPSYS_UNCONNECTED_124, SYNOPSYS_UNCONNECTED_125,
         SYNOPSYS_UNCONNECTED_126, SYNOPSYS_UNCONNECTED_127,
         SYNOPSYS_UNCONNECTED_128, SYNOPSYS_UNCONNECTED_129,
         SYNOPSYS_UNCONNECTED_130, SYNOPSYS_UNCONNECTED_131,
         SYNOPSYS_UNCONNECTED_132, SYNOPSYS_UNCONNECTED_133,
         SYNOPSYS_UNCONNECTED_134, SYNOPSYS_UNCONNECTED_135,
         SYNOPSYS_UNCONNECTED_136, SYNOPSYS_UNCONNECTED_137,
         SYNOPSYS_UNCONNECTED_138, SYNOPSYS_UNCONNECTED_139,
         SYNOPSYS_UNCONNECTED_140, SYNOPSYS_UNCONNECTED_141,
         SYNOPSYS_UNCONNECTED_142, SYNOPSYS_UNCONNECTED_143,
         SYNOPSYS_UNCONNECTED_144, SYNOPSYS_UNCONNECTED_145,
         SYNOPSYS_UNCONNECTED_146, SYNOPSYS_UNCONNECTED_147,
         SYNOPSYS_UNCONNECTED_148, SYNOPSYS_UNCONNECTED_149,
         SYNOPSYS_UNCONNECTED_150, SYNOPSYS_UNCONNECTED_151,
         SYNOPSYS_UNCONNECTED_152, SYNOPSYS_UNCONNECTED_153,
         SYNOPSYS_UNCONNECTED_154, SYNOPSYS_UNCONNECTED_155,
         SYNOPSYS_UNCONNECTED_156, SYNOPSYS_UNCONNECTED_157,
         SYNOPSYS_UNCONNECTED_158, SYNOPSYS_UNCONNECTED_159,
         SYNOPSYS_UNCONNECTED_160, SYNOPSYS_UNCONNECTED_161,
         SYNOPSYS_UNCONNECTED_162, SYNOPSYS_UNCONNECTED_163,
         SYNOPSYS_UNCONNECTED_164, SYNOPSYS_UNCONNECTED_165,
         SYNOPSYS_UNCONNECTED_166, SYNOPSYS_UNCONNECTED_167,
         SYNOPSYS_UNCONNECTED_168, SYNOPSYS_UNCONNECTED_169,
         SYNOPSYS_UNCONNECTED_170, SYNOPSYS_UNCONNECTED_171,
         SYNOPSYS_UNCONNECTED_172, SYNOPSYS_UNCONNECTED_173,
         SYNOPSYS_UNCONNECTED_174, SYNOPSYS_UNCONNECTED_175,
         SYNOPSYS_UNCONNECTED_176, SYNOPSYS_UNCONNECTED_177,
         SYNOPSYS_UNCONNECTED_178, SYNOPSYS_UNCONNECTED_179,
         SYNOPSYS_UNCONNECTED_180, SYNOPSYS_UNCONNECTED_181,
         SYNOPSYS_UNCONNECTED_182, SYNOPSYS_UNCONNECTED_183,
         SYNOPSYS_UNCONNECTED_184, SYNOPSYS_UNCONNECTED_185,
         SYNOPSYS_UNCONNECTED_186, SYNOPSYS_UNCONNECTED_187,
         SYNOPSYS_UNCONNECTED_188, SYNOPSYS_UNCONNECTED_189,
         SYNOPSYS_UNCONNECTED_190, SYNOPSYS_UNCONNECTED_191,
         SYNOPSYS_UNCONNECTED_192, SYNOPSYS_UNCONNECTED_193,
         SYNOPSYS_UNCONNECTED_194, SYNOPSYS_UNCONNECTED_195,
         SYNOPSYS_UNCONNECTED_196, SYNOPSYS_UNCONNECTED_197,
         SYNOPSYS_UNCONNECTED_198, SYNOPSYS_UNCONNECTED_199,
         SYNOPSYS_UNCONNECTED_200, SYNOPSYS_UNCONNECTED_201,
         SYNOPSYS_UNCONNECTED_202, SYNOPSYS_UNCONNECTED_203,
         SYNOPSYS_UNCONNECTED_204, SYNOPSYS_UNCONNECTED_205,
         SYNOPSYS_UNCONNECTED_206, SYNOPSYS_UNCONNECTED_207,
         SYNOPSYS_UNCONNECTED_208, SYNOPSYS_UNCONNECTED_209,
         SYNOPSYS_UNCONNECTED_210, SYNOPSYS_UNCONNECTED_211,
         SYNOPSYS_UNCONNECTED_212, SYNOPSYS_UNCONNECTED_213,
         SYNOPSYS_UNCONNECTED_214, SYNOPSYS_UNCONNECTED_215,
         SYNOPSYS_UNCONNECTED_216, SYNOPSYS_UNCONNECTED_217,
         SYNOPSYS_UNCONNECTED_218, SYNOPSYS_UNCONNECTED_219,
         SYNOPSYS_UNCONNECTED_220, SYNOPSYS_UNCONNECTED_221,
         SYNOPSYS_UNCONNECTED_222, SYNOPSYS_UNCONNECTED_223,
         SYNOPSYS_UNCONNECTED_224, SYNOPSYS_UNCONNECTED_225,
         SYNOPSYS_UNCONNECTED_226, SYNOPSYS_UNCONNECTED_227,
         SYNOPSYS_UNCONNECTED_228, SYNOPSYS_UNCONNECTED_229,
         SYNOPSYS_UNCONNECTED_230, SYNOPSYS_UNCONNECTED_231,
         SYNOPSYS_UNCONNECTED_232, SYNOPSYS_UNCONNECTED_233,
         SYNOPSYS_UNCONNECTED_234, SYNOPSYS_UNCONNECTED_235,
         SYNOPSYS_UNCONNECTED_236, SYNOPSYS_UNCONNECTED_237,
         SYNOPSYS_UNCONNECTED_238, SYNOPSYS_UNCONNECTED_239,
         SYNOPSYS_UNCONNECTED_240, SYNOPSYS_UNCONNECTED_241,
         SYNOPSYS_UNCONNECTED_242, SYNOPSYS_UNCONNECTED_243,
         SYNOPSYS_UNCONNECTED_244, SYNOPSYS_UNCONNECTED_245,
         SYNOPSYS_UNCONNECTED_246, SYNOPSYS_UNCONNECTED_247,
         SYNOPSYS_UNCONNECTED_248, SYNOPSYS_UNCONNECTED_249,
         SYNOPSYS_UNCONNECTED_250, SYNOPSYS_UNCONNECTED_251,
         SYNOPSYS_UNCONNECTED_252, SYNOPSYS_UNCONNECTED_253,
         SYNOPSYS_UNCONNECTED_254, SYNOPSYS_UNCONNECTED_255,
         SYNOPSYS_UNCONNECTED_256, SYNOPSYS_UNCONNECTED_257,
         SYNOPSYS_UNCONNECTED_258, SYNOPSYS_UNCONNECTED_259,
         SYNOPSYS_UNCONNECTED_260, SYNOPSYS_UNCONNECTED_261,
         SYNOPSYS_UNCONNECTED_262, SYNOPSYS_UNCONNECTED_263,
         SYNOPSYS_UNCONNECTED_264, SYNOPSYS_UNCONNECTED_265,
         SYNOPSYS_UNCONNECTED_266, SYNOPSYS_UNCONNECTED_267,
         SYNOPSYS_UNCONNECTED_268, SYNOPSYS_UNCONNECTED_269,
         SYNOPSYS_UNCONNECTED_270, SYNOPSYS_UNCONNECTED_271,
         SYNOPSYS_UNCONNECTED_272, SYNOPSYS_UNCONNECTED_273,
         SYNOPSYS_UNCONNECTED_274, SYNOPSYS_UNCONNECTED_275,
         SYNOPSYS_UNCONNECTED_276, SYNOPSYS_UNCONNECTED_277,
         SYNOPSYS_UNCONNECTED_278, SYNOPSYS_UNCONNECTED_279,
         SYNOPSYS_UNCONNECTED_280, SYNOPSYS_UNCONNECTED_281,
         SYNOPSYS_UNCONNECTED_282, SYNOPSYS_UNCONNECTED_283,
         SYNOPSYS_UNCONNECTED_284, SYNOPSYS_UNCONNECTED_285,
         SYNOPSYS_UNCONNECTED_286, SYNOPSYS_UNCONNECTED_287,
         SYNOPSYS_UNCONNECTED_288, SYNOPSYS_UNCONNECTED_289,
         SYNOPSYS_UNCONNECTED_290, SYNOPSYS_UNCONNECTED_291,
         SYNOPSYS_UNCONNECTED_292, SYNOPSYS_UNCONNECTED_293,
         SYNOPSYS_UNCONNECTED_294, SYNOPSYS_UNCONNECTED_295,
         SYNOPSYS_UNCONNECTED_296, SYNOPSYS_UNCONNECTED_297,
         SYNOPSYS_UNCONNECTED_298, SYNOPSYS_UNCONNECTED_299,
         SYNOPSYS_UNCONNECTED_300, SYNOPSYS_UNCONNECTED_301,
         SYNOPSYS_UNCONNECTED_302, SYNOPSYS_UNCONNECTED_303,
         SYNOPSYS_UNCONNECTED_304, SYNOPSYS_UNCONNECTED_305,
         SYNOPSYS_UNCONNECTED_306, SYNOPSYS_UNCONNECTED_307,
         SYNOPSYS_UNCONNECTED_308, SYNOPSYS_UNCONNECTED_309,
         SYNOPSYS_UNCONNECTED_310, SYNOPSYS_UNCONNECTED_311,
         SYNOPSYS_UNCONNECTED_312, SYNOPSYS_UNCONNECTED_313,
         SYNOPSYS_UNCONNECTED_314, SYNOPSYS_UNCONNECTED_315,
         SYNOPSYS_UNCONNECTED_316, SYNOPSYS_UNCONNECTED_317,
         SYNOPSYS_UNCONNECTED_318, SYNOPSYS_UNCONNECTED_319,
         SYNOPSYS_UNCONNECTED_320, SYNOPSYS_UNCONNECTED_321,
         SYNOPSYS_UNCONNECTED_322, SYNOPSYS_UNCONNECTED_323,
         SYNOPSYS_UNCONNECTED_324, SYNOPSYS_UNCONNECTED_325,
         SYNOPSYS_UNCONNECTED_326, SYNOPSYS_UNCONNECTED_327,
         SYNOPSYS_UNCONNECTED_328, SYNOPSYS_UNCONNECTED_329,
         SYNOPSYS_UNCONNECTED_330, SYNOPSYS_UNCONNECTED_331,
         SYNOPSYS_UNCONNECTED_332, SYNOPSYS_UNCONNECTED_333,
         SYNOPSYS_UNCONNECTED_334, SYNOPSYS_UNCONNECTED_335,
         SYNOPSYS_UNCONNECTED_336, SYNOPSYS_UNCONNECTED_337,
         SYNOPSYS_UNCONNECTED_338, SYNOPSYS_UNCONNECTED_339,
         SYNOPSYS_UNCONNECTED_340, SYNOPSYS_UNCONNECTED_341,
         SYNOPSYS_UNCONNECTED_342, SYNOPSYS_UNCONNECTED_343,
         SYNOPSYS_UNCONNECTED_344, SYNOPSYS_UNCONNECTED_345,
         SYNOPSYS_UNCONNECTED_346, SYNOPSYS_UNCONNECTED_347,
         SYNOPSYS_UNCONNECTED_348, SYNOPSYS_UNCONNECTED_349,
         SYNOPSYS_UNCONNECTED_350, SYNOPSYS_UNCONNECTED_351,
         SYNOPSYS_UNCONNECTED_352, SYNOPSYS_UNCONNECTED_353,
         SYNOPSYS_UNCONNECTED_354, SYNOPSYS_UNCONNECTED_355,
         SYNOPSYS_UNCONNECTED_356, SYNOPSYS_UNCONNECTED_357,
         SYNOPSYS_UNCONNECTED_358, SYNOPSYS_UNCONNECTED_359,
         SYNOPSYS_UNCONNECTED_360, SYNOPSYS_UNCONNECTED_361,
         SYNOPSYS_UNCONNECTED_362, SYNOPSYS_UNCONNECTED_363,
         SYNOPSYS_UNCONNECTED_364, SYNOPSYS_UNCONNECTED_365,
         SYNOPSYS_UNCONNECTED_366, SYNOPSYS_UNCONNECTED_367,
         SYNOPSYS_UNCONNECTED_368, SYNOPSYS_UNCONNECTED_369,
         SYNOPSYS_UNCONNECTED_370, SYNOPSYS_UNCONNECTED_371,
         SYNOPSYS_UNCONNECTED_372, SYNOPSYS_UNCONNECTED_373,
         SYNOPSYS_UNCONNECTED_374, SYNOPSYS_UNCONNECTED_375,
         SYNOPSYS_UNCONNECTED_376, SYNOPSYS_UNCONNECTED_377,
         SYNOPSYS_UNCONNECTED_378, SYNOPSYS_UNCONNECTED_379,
         SYNOPSYS_UNCONNECTED_380, SYNOPSYS_UNCONNECTED_381,
         SYNOPSYS_UNCONNECTED_382, SYNOPSYS_UNCONNECTED_383,
         SYNOPSYS_UNCONNECTED_384, SYNOPSYS_UNCONNECTED_385,
         SYNOPSYS_UNCONNECTED_386, SYNOPSYS_UNCONNECTED_387,
         SYNOPSYS_UNCONNECTED_388, SYNOPSYS_UNCONNECTED_389,
         SYNOPSYS_UNCONNECTED_390, SYNOPSYS_UNCONNECTED_391,
         SYNOPSYS_UNCONNECTED_392, SYNOPSYS_UNCONNECTED_393,
         SYNOPSYS_UNCONNECTED_394, SYNOPSYS_UNCONNECTED_395,
         SYNOPSYS_UNCONNECTED_396, SYNOPSYS_UNCONNECTED_397,
         SYNOPSYS_UNCONNECTED_398, SYNOPSYS_UNCONNECTED_399,
         SYNOPSYS_UNCONNECTED_400, SYNOPSYS_UNCONNECTED_401,
         SYNOPSYS_UNCONNECTED_402, SYNOPSYS_UNCONNECTED_403,
         SYNOPSYS_UNCONNECTED_404, SYNOPSYS_UNCONNECTED_405,
         SYNOPSYS_UNCONNECTED_406, SYNOPSYS_UNCONNECTED_407,
         SYNOPSYS_UNCONNECTED_408, SYNOPSYS_UNCONNECTED_409,
         SYNOPSYS_UNCONNECTED_410, SYNOPSYS_UNCONNECTED_411,
         SYNOPSYS_UNCONNECTED_412, SYNOPSYS_UNCONNECTED_413,
         SYNOPSYS_UNCONNECTED_414, SYNOPSYS_UNCONNECTED_415,
         SYNOPSYS_UNCONNECTED_416, SYNOPSYS_UNCONNECTED_417,
         SYNOPSYS_UNCONNECTED_418, SYNOPSYS_UNCONNECTED_419,
         SYNOPSYS_UNCONNECTED_420, SYNOPSYS_UNCONNECTED_421,
         SYNOPSYS_UNCONNECTED_422, SYNOPSYS_UNCONNECTED_423,
         SYNOPSYS_UNCONNECTED_424, SYNOPSYS_UNCONNECTED_425,
         SYNOPSYS_UNCONNECTED_426, SYNOPSYS_UNCONNECTED_427,
         SYNOPSYS_UNCONNECTED_428, SYNOPSYS_UNCONNECTED_429,
         SYNOPSYS_UNCONNECTED_430, SYNOPSYS_UNCONNECTED_431,
         SYNOPSYS_UNCONNECTED_432, SYNOPSYS_UNCONNECTED_433,
         SYNOPSYS_UNCONNECTED_434, SYNOPSYS_UNCONNECTED_435,
         SYNOPSYS_UNCONNECTED_436, SYNOPSYS_UNCONNECTED_437,
         SYNOPSYS_UNCONNECTED_438, SYNOPSYS_UNCONNECTED_439,
         SYNOPSYS_UNCONNECTED_440, SYNOPSYS_UNCONNECTED_441,
         SYNOPSYS_UNCONNECTED_442, SYNOPSYS_UNCONNECTED_443,
         SYNOPSYS_UNCONNECTED_444, SYNOPSYS_UNCONNECTED_445,
         SYNOPSYS_UNCONNECTED_446, SYNOPSYS_UNCONNECTED_447,
         SYNOPSYS_UNCONNECTED_448, SYNOPSYS_UNCONNECTED_449,
         SYNOPSYS_UNCONNECTED_450, SYNOPSYS_UNCONNECTED_451,
         SYNOPSYS_UNCONNECTED_452, SYNOPSYS_UNCONNECTED_453,
         SYNOPSYS_UNCONNECTED_454, SYNOPSYS_UNCONNECTED_455,
         SYNOPSYS_UNCONNECTED_456, SYNOPSYS_UNCONNECTED_457,
         SYNOPSYS_UNCONNECTED_458, SYNOPSYS_UNCONNECTED_459,
         SYNOPSYS_UNCONNECTED_460, SYNOPSYS_UNCONNECTED_461,
         SYNOPSYS_UNCONNECTED_462, SYNOPSYS_UNCONNECTED_463,
         SYNOPSYS_UNCONNECTED_464, SYNOPSYS_UNCONNECTED_465,
         SYNOPSYS_UNCONNECTED_466, SYNOPSYS_UNCONNECTED_467,
         SYNOPSYS_UNCONNECTED_468, SYNOPSYS_UNCONNECTED_469,
         SYNOPSYS_UNCONNECTED_470, SYNOPSYS_UNCONNECTED_471,
         SYNOPSYS_UNCONNECTED_472, SYNOPSYS_UNCONNECTED_473,
         SYNOPSYS_UNCONNECTED_474, SYNOPSYS_UNCONNECTED_475,
         SYNOPSYS_UNCONNECTED_476, SYNOPSYS_UNCONNECTED_477,
         SYNOPSYS_UNCONNECTED_478, SYNOPSYS_UNCONNECTED_479,
         SYNOPSYS_UNCONNECTED_480, SYNOPSYS_UNCONNECTED_481,
         SYNOPSYS_UNCONNECTED_482, SYNOPSYS_UNCONNECTED_483,
         SYNOPSYS_UNCONNECTED_484, SYNOPSYS_UNCONNECTED_485,
         SYNOPSYS_UNCONNECTED_486, SYNOPSYS_UNCONNECTED_487,
         SYNOPSYS_UNCONNECTED_488, SYNOPSYS_UNCONNECTED_489,
         SYNOPSYS_UNCONNECTED_490, SYNOPSYS_UNCONNECTED_491,
         SYNOPSYS_UNCONNECTED_492, SYNOPSYS_UNCONNECTED_493,
         SYNOPSYS_UNCONNECTED_494, SYNOPSYS_UNCONNECTED_495,
         SYNOPSYS_UNCONNECTED_496, SYNOPSYS_UNCONNECTED_497,
         SYNOPSYS_UNCONNECTED_498, SYNOPSYS_UNCONNECTED_499,
         SYNOPSYS_UNCONNECTED_500, SYNOPSYS_UNCONNECTED_501,
         SYNOPSYS_UNCONNECTED_502, SYNOPSYS_UNCONNECTED_503,
         SYNOPSYS_UNCONNECTED_504, SYNOPSYS_UNCONNECTED_505,
         SYNOPSYS_UNCONNECTED_506, SYNOPSYS_UNCONNECTED_507,
         SYNOPSYS_UNCONNECTED_508, SYNOPSYS_UNCONNECTED_509,
         SYNOPSYS_UNCONNECTED_510, SYNOPSYS_UNCONNECTED_511,
         SYNOPSYS_UNCONNECTED_512, SYNOPSYS_UNCONNECTED_513,
         SYNOPSYS_UNCONNECTED_514, SYNOPSYS_UNCONNECTED_515,
         SYNOPSYS_UNCONNECTED_516, SYNOPSYS_UNCONNECTED_517,
         SYNOPSYS_UNCONNECTED_518, SYNOPSYS_UNCONNECTED_519,
         SYNOPSYS_UNCONNECTED_520, SYNOPSYS_UNCONNECTED_521,
         SYNOPSYS_UNCONNECTED_522, SYNOPSYS_UNCONNECTED_523,
         SYNOPSYS_UNCONNECTED_524, SYNOPSYS_UNCONNECTED_525,
         SYNOPSYS_UNCONNECTED_526, SYNOPSYS_UNCONNECTED_527,
         SYNOPSYS_UNCONNECTED_528, SYNOPSYS_UNCONNECTED_529,
         SYNOPSYS_UNCONNECTED_530, SYNOPSYS_UNCONNECTED_531,
         SYNOPSYS_UNCONNECTED_532, SYNOPSYS_UNCONNECTED_533,
         SYNOPSYS_UNCONNECTED_534, SYNOPSYS_UNCONNECTED_535,
         SYNOPSYS_UNCONNECTED_536, SYNOPSYS_UNCONNECTED_537,
         SYNOPSYS_UNCONNECTED_538, SYNOPSYS_UNCONNECTED_539,
         SYNOPSYS_UNCONNECTED_540, SYNOPSYS_UNCONNECTED_541,
         SYNOPSYS_UNCONNECTED_542, SYNOPSYS_UNCONNECTED_543,
         SYNOPSYS_UNCONNECTED_544, SYNOPSYS_UNCONNECTED_545,
         SYNOPSYS_UNCONNECTED_546, SYNOPSYS_UNCONNECTED_547,
         SYNOPSYS_UNCONNECTED_548, SYNOPSYS_UNCONNECTED_549,
         SYNOPSYS_UNCONNECTED_550, SYNOPSYS_UNCONNECTED_551,
         SYNOPSYS_UNCONNECTED_552, SYNOPSYS_UNCONNECTED_553,
         SYNOPSYS_UNCONNECTED_554, SYNOPSYS_UNCONNECTED_555,
         SYNOPSYS_UNCONNECTED_556, SYNOPSYS_UNCONNECTED_557,
         SYNOPSYS_UNCONNECTED_558, SYNOPSYS_UNCONNECTED_559,
         SYNOPSYS_UNCONNECTED_560, SYNOPSYS_UNCONNECTED_561,
         SYNOPSYS_UNCONNECTED_562, SYNOPSYS_UNCONNECTED_563,
         SYNOPSYS_UNCONNECTED_564, SYNOPSYS_UNCONNECTED_565,
         SYNOPSYS_UNCONNECTED_566, SYNOPSYS_UNCONNECTED_567,
         SYNOPSYS_UNCONNECTED_568, SYNOPSYS_UNCONNECTED_569,
         SYNOPSYS_UNCONNECTED_570, SYNOPSYS_UNCONNECTED_571,
         SYNOPSYS_UNCONNECTED_572, SYNOPSYS_UNCONNECTED_573,
         SYNOPSYS_UNCONNECTED_574, SYNOPSYS_UNCONNECTED_575,
         SYNOPSYS_UNCONNECTED_576, SYNOPSYS_UNCONNECTED_577,
         SYNOPSYS_UNCONNECTED_578, SYNOPSYS_UNCONNECTED_579,
         SYNOPSYS_UNCONNECTED_580, SYNOPSYS_UNCONNECTED_581,
         SYNOPSYS_UNCONNECTED_582, SYNOPSYS_UNCONNECTED_583,
         SYNOPSYS_UNCONNECTED_584, SYNOPSYS_UNCONNECTED_585,
         SYNOPSYS_UNCONNECTED_586, SYNOPSYS_UNCONNECTED_587,
         SYNOPSYS_UNCONNECTED_588, SYNOPSYS_UNCONNECTED_589,
         SYNOPSYS_UNCONNECTED_590, SYNOPSYS_UNCONNECTED_591,
         SYNOPSYS_UNCONNECTED_592, SYNOPSYS_UNCONNECTED_593,
         SYNOPSYS_UNCONNECTED_594, SYNOPSYS_UNCONNECTED_595,
         SYNOPSYS_UNCONNECTED_596, SYNOPSYS_UNCONNECTED_597,
         SYNOPSYS_UNCONNECTED_598, SYNOPSYS_UNCONNECTED_599,
         SYNOPSYS_UNCONNECTED_600, SYNOPSYS_UNCONNECTED_601,
         SYNOPSYS_UNCONNECTED_602, SYNOPSYS_UNCONNECTED_603,
         SYNOPSYS_UNCONNECTED_604, SYNOPSYS_UNCONNECTED_605,
         SYNOPSYS_UNCONNECTED_606, SYNOPSYS_UNCONNECTED_607,
         SYNOPSYS_UNCONNECTED_608, SYNOPSYS_UNCONNECTED_609,
         SYNOPSYS_UNCONNECTED_610, SYNOPSYS_UNCONNECTED_611,
         SYNOPSYS_UNCONNECTED_612, SYNOPSYS_UNCONNECTED_613,
         SYNOPSYS_UNCONNECTED_614, SYNOPSYS_UNCONNECTED_615,
         SYNOPSYS_UNCONNECTED_616, SYNOPSYS_UNCONNECTED_617,
         SYNOPSYS_UNCONNECTED_618, SYNOPSYS_UNCONNECTED_619,
         SYNOPSYS_UNCONNECTED_620, SYNOPSYS_UNCONNECTED_621,
         SYNOPSYS_UNCONNECTED_622, SYNOPSYS_UNCONNECTED_623,
         SYNOPSYS_UNCONNECTED_624, SYNOPSYS_UNCONNECTED_625,
         SYNOPSYS_UNCONNECTED_626, SYNOPSYS_UNCONNECTED_627,
         SYNOPSYS_UNCONNECTED_628, SYNOPSYS_UNCONNECTED_629,
         SYNOPSYS_UNCONNECTED_630, SYNOPSYS_UNCONNECTED_631,
         SYNOPSYS_UNCONNECTED_632, SYNOPSYS_UNCONNECTED_633,
         SYNOPSYS_UNCONNECTED_634, SYNOPSYS_UNCONNECTED_635,
         SYNOPSYS_UNCONNECTED_636, SYNOPSYS_UNCONNECTED_637,
         SYNOPSYS_UNCONNECTED_638, SYNOPSYS_UNCONNECTED_639,
         SYNOPSYS_UNCONNECTED_640, SYNOPSYS_UNCONNECTED_641,
         SYNOPSYS_UNCONNECTED_642, SYNOPSYS_UNCONNECTED_643,
         SYNOPSYS_UNCONNECTED_644, SYNOPSYS_UNCONNECTED_645,
         SYNOPSYS_UNCONNECTED_646, SYNOPSYS_UNCONNECTED_647,
         SYNOPSYS_UNCONNECTED_648, SYNOPSYS_UNCONNECTED_649,
         SYNOPSYS_UNCONNECTED_650, SYNOPSYS_UNCONNECTED_651,
         SYNOPSYS_UNCONNECTED_652, SYNOPSYS_UNCONNECTED_653,
         SYNOPSYS_UNCONNECTED_654, SYNOPSYS_UNCONNECTED_655,
         SYNOPSYS_UNCONNECTED_656, SYNOPSYS_UNCONNECTED_657,
         SYNOPSYS_UNCONNECTED_658, SYNOPSYS_UNCONNECTED_659,
         SYNOPSYS_UNCONNECTED_660, SYNOPSYS_UNCONNECTED_661,
         SYNOPSYS_UNCONNECTED_662, SYNOPSYS_UNCONNECTED_663,
         SYNOPSYS_UNCONNECTED_664, SYNOPSYS_UNCONNECTED_665,
         SYNOPSYS_UNCONNECTED_666, SYNOPSYS_UNCONNECTED_667,
         SYNOPSYS_UNCONNECTED_668, SYNOPSYS_UNCONNECTED_669,
         SYNOPSYS_UNCONNECTED_670, SYNOPSYS_UNCONNECTED_671,
         SYNOPSYS_UNCONNECTED_672, SYNOPSYS_UNCONNECTED_673,
         SYNOPSYS_UNCONNECTED_674, SYNOPSYS_UNCONNECTED_675,
         SYNOPSYS_UNCONNECTED_676, SYNOPSYS_UNCONNECTED_677,
         SYNOPSYS_UNCONNECTED_678, SYNOPSYS_UNCONNECTED_679,
         SYNOPSYS_UNCONNECTED_680, SYNOPSYS_UNCONNECTED_681,
         SYNOPSYS_UNCONNECTED_682, SYNOPSYS_UNCONNECTED_683,
         SYNOPSYS_UNCONNECTED_684, SYNOPSYS_UNCONNECTED_685,
         SYNOPSYS_UNCONNECTED_686, SYNOPSYS_UNCONNECTED_687,
         SYNOPSYS_UNCONNECTED_688, SYNOPSYS_UNCONNECTED_689,
         SYNOPSYS_UNCONNECTED_690, SYNOPSYS_UNCONNECTED_691,
         SYNOPSYS_UNCONNECTED_692, SYNOPSYS_UNCONNECTED_693,
         SYNOPSYS_UNCONNECTED_694, SYNOPSYS_UNCONNECTED_695,
         SYNOPSYS_UNCONNECTED_696, SYNOPSYS_UNCONNECTED_697,
         SYNOPSYS_UNCONNECTED_698, SYNOPSYS_UNCONNECTED_699,
         SYNOPSYS_UNCONNECTED_700, SYNOPSYS_UNCONNECTED_701,
         SYNOPSYS_UNCONNECTED_702, SYNOPSYS_UNCONNECTED_703,
         SYNOPSYS_UNCONNECTED_704, SYNOPSYS_UNCONNECTED_705,
         SYNOPSYS_UNCONNECTED_706, SYNOPSYS_UNCONNECTED_707,
         SYNOPSYS_UNCONNECTED_708, SYNOPSYS_UNCONNECTED_709,
         SYNOPSYS_UNCONNECTED_710, SYNOPSYS_UNCONNECTED_711,
         SYNOPSYS_UNCONNECTED_712, SYNOPSYS_UNCONNECTED_713,
         SYNOPSYS_UNCONNECTED_714, SYNOPSYS_UNCONNECTED_715,
         SYNOPSYS_UNCONNECTED_716, SYNOPSYS_UNCONNECTED_717,
         SYNOPSYS_UNCONNECTED_718, SYNOPSYS_UNCONNECTED_719,
         SYNOPSYS_UNCONNECTED_720, SYNOPSYS_UNCONNECTED_721,
         SYNOPSYS_UNCONNECTED_722, SYNOPSYS_UNCONNECTED_723,
         SYNOPSYS_UNCONNECTED_724, SYNOPSYS_UNCONNECTED_725,
         SYNOPSYS_UNCONNECTED_726, SYNOPSYS_UNCONNECTED_727,
         SYNOPSYS_UNCONNECTED_728, SYNOPSYS_UNCONNECTED_729,
         SYNOPSYS_UNCONNECTED_730, SYNOPSYS_UNCONNECTED_731,
         SYNOPSYS_UNCONNECTED_732, SYNOPSYS_UNCONNECTED_733,
         SYNOPSYS_UNCONNECTED_734, SYNOPSYS_UNCONNECTED_735,
         SYNOPSYS_UNCONNECTED_736, SYNOPSYS_UNCONNECTED_737,
         SYNOPSYS_UNCONNECTED_738, SYNOPSYS_UNCONNECTED_739,
         SYNOPSYS_UNCONNECTED_740, SYNOPSYS_UNCONNECTED_741,
         SYNOPSYS_UNCONNECTED_742, SYNOPSYS_UNCONNECTED_743,
         SYNOPSYS_UNCONNECTED_744, SYNOPSYS_UNCONNECTED_745,
         SYNOPSYS_UNCONNECTED_746, SYNOPSYS_UNCONNECTED_747,
         SYNOPSYS_UNCONNECTED_748, SYNOPSYS_UNCONNECTED_749,
         SYNOPSYS_UNCONNECTED_750, SYNOPSYS_UNCONNECTED_751,
         SYNOPSYS_UNCONNECTED_752, SYNOPSYS_UNCONNECTED_753,
         SYNOPSYS_UNCONNECTED_754, SYNOPSYS_UNCONNECTED_755,
         SYNOPSYS_UNCONNECTED_756, SYNOPSYS_UNCONNECTED_757,
         SYNOPSYS_UNCONNECTED_758, SYNOPSYS_UNCONNECTED_759,
         SYNOPSYS_UNCONNECTED_760, SYNOPSYS_UNCONNECTED_761,
         SYNOPSYS_UNCONNECTED_762, SYNOPSYS_UNCONNECTED_763,
         SYNOPSYS_UNCONNECTED_764, SYNOPSYS_UNCONNECTED_765,
         SYNOPSYS_UNCONNECTED_766, SYNOPSYS_UNCONNECTED_767,
         SYNOPSYS_UNCONNECTED_768, SYNOPSYS_UNCONNECTED_769,
         SYNOPSYS_UNCONNECTED_770, SYNOPSYS_UNCONNECTED_771,
         SYNOPSYS_UNCONNECTED_772, SYNOPSYS_UNCONNECTED_773,
         SYNOPSYS_UNCONNECTED_774, SYNOPSYS_UNCONNECTED_775,
         SYNOPSYS_UNCONNECTED_776, SYNOPSYS_UNCONNECTED_777,
         SYNOPSYS_UNCONNECTED_778, SYNOPSYS_UNCONNECTED_779,
         SYNOPSYS_UNCONNECTED_780, SYNOPSYS_UNCONNECTED_781,
         SYNOPSYS_UNCONNECTED_782, SYNOPSYS_UNCONNECTED_783,
         SYNOPSYS_UNCONNECTED_784, SYNOPSYS_UNCONNECTED_785,
         SYNOPSYS_UNCONNECTED_786, SYNOPSYS_UNCONNECTED_787,
         SYNOPSYS_UNCONNECTED_788, SYNOPSYS_UNCONNECTED_789,
         SYNOPSYS_UNCONNECTED_790, SYNOPSYS_UNCONNECTED_791,
         SYNOPSYS_UNCONNECTED_792, SYNOPSYS_UNCONNECTED_793,
         SYNOPSYS_UNCONNECTED_794, SYNOPSYS_UNCONNECTED_795,
         SYNOPSYS_UNCONNECTED_796, SYNOPSYS_UNCONNECTED_797,
         SYNOPSYS_UNCONNECTED_798, SYNOPSYS_UNCONNECTED_799,
         SYNOPSYS_UNCONNECTED_800, SYNOPSYS_UNCONNECTED_801,
         SYNOPSYS_UNCONNECTED_802, SYNOPSYS_UNCONNECTED_803,
         SYNOPSYS_UNCONNECTED_804, SYNOPSYS_UNCONNECTED_805,
         SYNOPSYS_UNCONNECTED_806, SYNOPSYS_UNCONNECTED_807,
         SYNOPSYS_UNCONNECTED_808, SYNOPSYS_UNCONNECTED_809,
         SYNOPSYS_UNCONNECTED_810, SYNOPSYS_UNCONNECTED_811,
         SYNOPSYS_UNCONNECTED_812, SYNOPSYS_UNCONNECTED_813,
         SYNOPSYS_UNCONNECTED_814, SYNOPSYS_UNCONNECTED_815,
         SYNOPSYS_UNCONNECTED_816, SYNOPSYS_UNCONNECTED_817,
         SYNOPSYS_UNCONNECTED_818, SYNOPSYS_UNCONNECTED_819,
         SYNOPSYS_UNCONNECTED_820, SYNOPSYS_UNCONNECTED_821,
         SYNOPSYS_UNCONNECTED_822, SYNOPSYS_UNCONNECTED_823,
         SYNOPSYS_UNCONNECTED_824, SYNOPSYS_UNCONNECTED_825,
         SYNOPSYS_UNCONNECTED_826, SYNOPSYS_UNCONNECTED_827,
         SYNOPSYS_UNCONNECTED_828, SYNOPSYS_UNCONNECTED_829,
         SYNOPSYS_UNCONNECTED_830, SYNOPSYS_UNCONNECTED_831,
         SYNOPSYS_UNCONNECTED_832, SYNOPSYS_UNCONNECTED_833,
         SYNOPSYS_UNCONNECTED_834, SYNOPSYS_UNCONNECTED_835,
         SYNOPSYS_UNCONNECTED_836, SYNOPSYS_UNCONNECTED_837,
         SYNOPSYS_UNCONNECTED_838, SYNOPSYS_UNCONNECTED_839,
         SYNOPSYS_UNCONNECTED_840, SYNOPSYS_UNCONNECTED_841,
         SYNOPSYS_UNCONNECTED_842, SYNOPSYS_UNCONNECTED_843,
         SYNOPSYS_UNCONNECTED_844, SYNOPSYS_UNCONNECTED_845,
         SYNOPSYS_UNCONNECTED_846, SYNOPSYS_UNCONNECTED_847,
         SYNOPSYS_UNCONNECTED_848, SYNOPSYS_UNCONNECTED_849,
         SYNOPSYS_UNCONNECTED_850, SYNOPSYS_UNCONNECTED_851,
         SYNOPSYS_UNCONNECTED_852, SYNOPSYS_UNCONNECTED_853,
         SYNOPSYS_UNCONNECTED_854, SYNOPSYS_UNCONNECTED_855,
         SYNOPSYS_UNCONNECTED_856, SYNOPSYS_UNCONNECTED_857,
         SYNOPSYS_UNCONNECTED_858, SYNOPSYS_UNCONNECTED_859,
         SYNOPSYS_UNCONNECTED_860, SYNOPSYS_UNCONNECTED_861,
         SYNOPSYS_UNCONNECTED_862, SYNOPSYS_UNCONNECTED_863,
         SYNOPSYS_UNCONNECTED_864, SYNOPSYS_UNCONNECTED_865,
         SYNOPSYS_UNCONNECTED_866, SYNOPSYS_UNCONNECTED_867,
         SYNOPSYS_UNCONNECTED_868, SYNOPSYS_UNCONNECTED_869,
         SYNOPSYS_UNCONNECTED_870, SYNOPSYS_UNCONNECTED_871,
         SYNOPSYS_UNCONNECTED_872, SYNOPSYS_UNCONNECTED_873,
         SYNOPSYS_UNCONNECTED_874, SYNOPSYS_UNCONNECTED_875,
         SYNOPSYS_UNCONNECTED_876, SYNOPSYS_UNCONNECTED_877,
         SYNOPSYS_UNCONNECTED_878, SYNOPSYS_UNCONNECTED_879,
         SYNOPSYS_UNCONNECTED_880, SYNOPSYS_UNCONNECTED_881,
         SYNOPSYS_UNCONNECTED_882, SYNOPSYS_UNCONNECTED_883,
         SYNOPSYS_UNCONNECTED_884, SYNOPSYS_UNCONNECTED_885,
         SYNOPSYS_UNCONNECTED_886, SYNOPSYS_UNCONNECTED_887,
         SYNOPSYS_UNCONNECTED_888, SYNOPSYS_UNCONNECTED_889,
         SYNOPSYS_UNCONNECTED_890, SYNOPSYS_UNCONNECTED_891,
         SYNOPSYS_UNCONNECTED_892, SYNOPSYS_UNCONNECTED_893,
         SYNOPSYS_UNCONNECTED_894, SYNOPSYS_UNCONNECTED_895,
         SYNOPSYS_UNCONNECTED_896, SYNOPSYS_UNCONNECTED_897,
         SYNOPSYS_UNCONNECTED_898, SYNOPSYS_UNCONNECTED_899,
         SYNOPSYS_UNCONNECTED_900, SYNOPSYS_UNCONNECTED_901,
         SYNOPSYS_UNCONNECTED_902, SYNOPSYS_UNCONNECTED_903,
         SYNOPSYS_UNCONNECTED_904, SYNOPSYS_UNCONNECTED_905,
         SYNOPSYS_UNCONNECTED_906, SYNOPSYS_UNCONNECTED_907,
         SYNOPSYS_UNCONNECTED_908, SYNOPSYS_UNCONNECTED_909,
         SYNOPSYS_UNCONNECTED_910, SYNOPSYS_UNCONNECTED_911,
         SYNOPSYS_UNCONNECTED_912, SYNOPSYS_UNCONNECTED_913,
         SYNOPSYS_UNCONNECTED_914, SYNOPSYS_UNCONNECTED_915,
         SYNOPSYS_UNCONNECTED_916, SYNOPSYS_UNCONNECTED_917,
         SYNOPSYS_UNCONNECTED_918, SYNOPSYS_UNCONNECTED_919,
         SYNOPSYS_UNCONNECTED_920, SYNOPSYS_UNCONNECTED_921,
         SYNOPSYS_UNCONNECTED_922, SYNOPSYS_UNCONNECTED_923,
         SYNOPSYS_UNCONNECTED_924, SYNOPSYS_UNCONNECTED_925,
         SYNOPSYS_UNCONNECTED_926, SYNOPSYS_UNCONNECTED_927,
         SYNOPSYS_UNCONNECTED_928, SYNOPSYS_UNCONNECTED_929,
         SYNOPSYS_UNCONNECTED_930, SYNOPSYS_UNCONNECTED_931,
         SYNOPSYS_UNCONNECTED_932, SYNOPSYS_UNCONNECTED_933,
         SYNOPSYS_UNCONNECTED_934, SYNOPSYS_UNCONNECTED_935,
         SYNOPSYS_UNCONNECTED_936, SYNOPSYS_UNCONNECTED_937,
         SYNOPSYS_UNCONNECTED_938, SYNOPSYS_UNCONNECTED_939,
         SYNOPSYS_UNCONNECTED_940, SYNOPSYS_UNCONNECTED_941,
         SYNOPSYS_UNCONNECTED_942, SYNOPSYS_UNCONNECTED_943,
         SYNOPSYS_UNCONNECTED_944, SYNOPSYS_UNCONNECTED_945,
         SYNOPSYS_UNCONNECTED_946, SYNOPSYS_UNCONNECTED_947,
         SYNOPSYS_UNCONNECTED_948, SYNOPSYS_UNCONNECTED_949,
         SYNOPSYS_UNCONNECTED_950, SYNOPSYS_UNCONNECTED_951,
         SYNOPSYS_UNCONNECTED_952, SYNOPSYS_UNCONNECTED_953,
         SYNOPSYS_UNCONNECTED_954, SYNOPSYS_UNCONNECTED_955,
         SYNOPSYS_UNCONNECTED_956, SYNOPSYS_UNCONNECTED_957,
         SYNOPSYS_UNCONNECTED_958, SYNOPSYS_UNCONNECTED_959,
         SYNOPSYS_UNCONNECTED_960, SYNOPSYS_UNCONNECTED_961,
         SYNOPSYS_UNCONNECTED_962, SYNOPSYS_UNCONNECTED_963,
         SYNOPSYS_UNCONNECTED_964, SYNOPSYS_UNCONNECTED_965,
         SYNOPSYS_UNCONNECTED_966, SYNOPSYS_UNCONNECTED_967,
         SYNOPSYS_UNCONNECTED_968, SYNOPSYS_UNCONNECTED_969,
         SYNOPSYS_UNCONNECTED_970, SYNOPSYS_UNCONNECTED_971,
         SYNOPSYS_UNCONNECTED_972, SYNOPSYS_UNCONNECTED_973,
         SYNOPSYS_UNCONNECTED_974, SYNOPSYS_UNCONNECTED_975,
         SYNOPSYS_UNCONNECTED_976, SYNOPSYS_UNCONNECTED_977,
         SYNOPSYS_UNCONNECTED_978, SYNOPSYS_UNCONNECTED_979,
         SYNOPSYS_UNCONNECTED_980, SYNOPSYS_UNCONNECTED_981,
         SYNOPSYS_UNCONNECTED_982, SYNOPSYS_UNCONNECTED_983,
         SYNOPSYS_UNCONNECTED_984, SYNOPSYS_UNCONNECTED_985,
         SYNOPSYS_UNCONNECTED_986, SYNOPSYS_UNCONNECTED_987,
         SYNOPSYS_UNCONNECTED_988, SYNOPSYS_UNCONNECTED_989,
         SYNOPSYS_UNCONNECTED_990, SYNOPSYS_UNCONNECTED_991,
         SYNOPSYS_UNCONNECTED_992, SYNOPSYS_UNCONNECTED_993,
         SYNOPSYS_UNCONNECTED_994, SYNOPSYS_UNCONNECTED_995,
         SYNOPSYS_UNCONNECTED_996, SYNOPSYS_UNCONNECTED_997,
         SYNOPSYS_UNCONNECTED_998, SYNOPSYS_UNCONNECTED_999,
         SYNOPSYS_UNCONNECTED_1000, SYNOPSYS_UNCONNECTED_1001,
         SYNOPSYS_UNCONNECTED_1002, SYNOPSYS_UNCONNECTED_1003,
         SYNOPSYS_UNCONNECTED_1004, SYNOPSYS_UNCONNECTED_1005,
         SYNOPSYS_UNCONNECTED_1006, SYNOPSYS_UNCONNECTED_1007,
         SYNOPSYS_UNCONNECTED_1008, SYNOPSYS_UNCONNECTED_1009,
         SYNOPSYS_UNCONNECTED_1010, SYNOPSYS_UNCONNECTED_1011,
         SYNOPSYS_UNCONNECTED_1012, SYNOPSYS_UNCONNECTED_1013,
         SYNOPSYS_UNCONNECTED_1014, SYNOPSYS_UNCONNECTED_1015,
         SYNOPSYS_UNCONNECTED_1016, SYNOPSYS_UNCONNECTED_1017;
  wire   [183:174] hit;
  wire   [167:162] we;
  wire   [3:2] regE3;
  wire   [7:0] regDF;
  wire   [7:0] regDE;
  wire   [7:0] regD4;
  wire   [7:0] reg31;
  wire   [7:0] reg30;
  wire   [7:0] reg28;
  wire   [7:0] reg27;
  wire   [7:1] reg21;
  wire   [4:0] reg20;
  wire   [7:3] reg12;
  wire   [7:0] reg06;
  wire   [7:0] reg05;
  wire   [7:0] regAF;
  wire   [7:0] regAE;
  wire   [5:0] regAD;
  wire   [7:0] regAC;
  wire   [7:0] regAB;
  wire   [7:0] reg94;
  wire   [7:0] irqAE;
  wire   [7:0] irqDF;
  wire   [7:0] irq28;
  wire   [7:0] irq04;
  wire   [7:0] irq03;
  wire   [1:0] drstz;
  wire   [4:0] rstcnt;
  wire   [1:0] r_phyrst;
  wire   [7:0] wd01;
  wire   [7:0] clr03;
  wire   [7:0] set03;
  wire   [7:0] clr04;
  wire   [7:0] set04;
  wire   [7:0] wd12;
  wire   [14:0] inst_ofs_plus;
  wire   [7:0] wd18;
  wire   [7:0] wd19;
  wire   [7:0] wd20;
  wire   [7:0] wd21;
  wire   [7:0] clr28;
  wire   [2:0] oscdwn_shft;
  wire   [3:0] osc_gate_n;
  wire   [7:0] d_p0;
  wire   [7:0] setDF;
  wire   [7:0] clrDF;
  wire   [7:0] clrAE;
  wire   [5:0] setAE;
  wire   [3:0] lt_regE4_3_0;
  wire   [4:2] add_179_carry;

  AND2X1 U0_MASK_0 ( .A(oscdwn_shft[2]), .B(as_p0_chg), .Y(p0_chg_clr) );
  AND2X1 U0_MASK_1 ( .A(regD4[7]), .B(di_stbovp), .Y(di_stbovp_clr) );
  AND2X1 U0_MASK_2 ( .A(regD4[6]), .B(di_rd_det), .Y(di_rd_det_clr) );
  AND2X1 U0_MASK_3 ( .A(r_srcctl[7]), .B(dmf_wkup), .Y(dm_fault_clr) );
  AND2X1 U0_MASK_4 ( .A(regD4[5]), .B(aswkup), .Y(osc_low_clr) );
  glreg_a0_79 u0_reg00 ( .clk(clk), .arstz(n103), .we(we_176), .wdat({n197, 
        n191, n188, n181, n174, n168, n163, n160}), .rdat({r_txendk, r_txauto}) );
  glreg_a0_78 u0_reg01 ( .clk(clk), .arstz(n85), .we(upd01), .wdat(wd01), 
        .rdat({r_last, r_first, r_unlock, r_txnumk}) );
  glsta_a0_6 u0_reg03 ( .clk(clk), .arstz(n92), .rst0(n16), .set2({set03[7:4], 
        n1120, set03[2:0]}), .clr1(clr03), .rdat(dbgpo[7:0]), .irq(irq03) );
  glsta_a0_5 u0_reg04 ( .clk(clk), .arstz(n86), .rst0(phyrst), .set2(set04), 
        .clr1(clr04), .rdat(dbgpo[15:8]), .irq(irq04) );
  glreg_a0_77 u0_reg05 ( .clk(clk), .arstz(n87), .we(we_181), .wdat({n197, 
        n191, n186, n180, n177, n168, sfr_wdat[1:0]}), .rdat(reg05) );
  glreg_a0_76 u0_reg06 ( .clk(clk), .arstz(n88), .we(we_182), .wdat({n197, 
        n191, n186, n180, n174, n168, sfr_wdat[1:0]}), .rdat(reg06) );
  glreg_a0_75 u0_reg11 ( .clk(clk), .arstz(n93), .we(we_187), .wdat({n197, 
        n191, n186, n180, n174, n168, sfr_wdat[1:0]}), .rdat({reg11_7_, 
        r_rxords_ena[6:5], reg11_4, r_rxords_ena[3:0]}) );
  glreg_a0_74 u0_reg12 ( .clk(clk), .arstz(n97), .we(upd12), .wdat(wd12), 
        .rdat({reg12, r_txshrt, reg12_1, r_pshords}) );
  glreg_WIDTH5_2 u0_reg14 ( .clk(clk), .arstz(n127), .we(r_set_cpmsgid), 
        .wdat({n197, n191, n186, n180, n174}), .rdat({r_auto_gdcrc[0], 
        r_auto_discard, r_spec, r_auto_gdcrc[1]}) );
  glreg_a0_73 u0_reg15 ( .clk(clk), .arstz(n99), .we(we_191), .wdat({n197, 
        n191, n186, n180, sfr_wdat[3], n168, sfr_wdat[1:0]}), .rdat(
        dbgpo[31:24]) );
  glreg_a0_72 u0_reg18 ( .clk(clk), .arstz(n100), .we(upd18), .wdat(wd18), 
        .rdat(r_inst_ofs[7:0]) );
  glreg_a0_71 u0_reg19 ( .clk(clk), .arstz(n101), .we(upd19), .wdat(wd19), 
        .rdat({reg19_7_, r_inst_ofs[14:8]}) );
  glreg_a0_70 u0_reg20 ( .clk(clk), .arstz(n106), .we(upd20), .wdat(wd20), 
        .rdat({r_dat_spec, r_dat_datarole, reg20}) );
  glreg_a0_69 u0_reg21 ( .clk(clk), .arstz(n112), .we(upd21), .wdat(wd21), 
        .rdat({reg21, r_dat_portrole}) );
  glreg_6_00000018 u0_reg25 ( .clk(clk), .arstz(n122), .we(n1096), .wdat({n186, 
        n183, n176, n168, n165, sfr_wdat[0]}), .rdat({r_i2c_attr, r_pg0_sel, 
        reg25_0_}) );
  glreg_WIDTH1_6 u0_reg26 ( .clk(clk), .arstz(n134), .we(n1095), .wdat(n160), 
        .rdat(lt_reg26_0) );
  glreg_1_1 u1_reg26 ( .clk(clk), .arstz(n134), .we(i2c_mode_upd), .wdat(
        i2c_mode_wdat), .rdat(r_hwi2c_en) );
  glreg_7_70 u2_reg26 ( .clk(clk), .arstz(n121), .we(n1095), .wdat({n200, n194, 
        n188, n180, n177, n168, n165}), .rdat(r_i2c_deva) );
  glreg_a0_68 u0_reg27 ( .clk(clk), .arstz(n120), .we(we_203), .wdat({n197, 
        n191, n186, n180, n177, n169, n165, n158}), .rdat(reg27) );
  glsta_a0_4 u0_reg28 ( .clk(clk), .arstz(n119), .rst0(1'b0), .set2(i2c_ev), 
        .clr1(clr28), .rdat(reg28), .irq(irq28) );
  glreg_a0_67 u0_reg31 ( .clk(clk), .arstz(n118), .we(upd31), .wdat(i_pc[15:8]), .rdat(reg31) );
  glreg_8_00000001 u0_regD1 ( .clk(clk), .arstz(n83), .we(we_209), .wdat({n197, 
        n191, n186, n180, n177, n169, n165, n160}), .rdat({r_exist1st, 
        r_ordrs4, r_strtch, r_bclk_sel, r_gpio_tm, r_gpio_oe[6], r_gpio_pu[6], 
        r_gpio_pd[6]}) );
  glreg_8_00000011 u0_regD3 ( .clk(clk), .arstz(n82), .we(we_211), .wdat({n197, 
        n191, n186, n183, n177, n169, n163, n160}), .rdat({regD3_7_, 
        r_gpio_oe[5], r_gpio_pu[5], r_gpio_pd[5], regD3_3, r_gpio_oe[4], 
        r_gpio_pu[4], r_gpio_pd[4]}) );
  glreg_WIDTH3 u4_regD4 ( .clk(clk), .arstz(n134), .we(n4), .wdat({n198, n192, 
        sfr_wdat[5]}), .rdat(regD4[7:5]) );
  glreg_WIDTH2_2 u3_regD4 ( .clk(clk), .arstz(pwrdn_rstz), .we(n4), .wdat({
        n180, n174}), .rdat(regD4[4:3]) );
  glreg_WIDTH1_5 u2_regD4 ( .clk(clk), .arstz(pwrdn_rstz), .we(n4), .wdat(n168), .rdat(regD4[2]) );
  glreg_WIDTH1_4 u1_regD4 ( .clk(clk), .arstz(osc_low_rstz), .we(n4), .wdat(
        n165), .rdat(regD4[1]) );
  glreg_WIDTH1_3 u0_regD4 ( .clk(clk), .arstz(pwrdn_rstz), .we(n4), .wdat(n160), .rdat(regD4[0]) );
  glreg_8_000000f0 u0_regD5 ( .clk(clk), .arstz(n78), .we(we_213), .wdat({n200, 
        n194, n188, n183, n177, n169, n163, n158}), .rdat({r_gpio_pu[3:0], 
        r_gpio_pd[3:0]}) );
  glreg_8_00000098 u0_regD6 ( .clk(clk), .arstz(n80), .we(we_214), .wdat({n200, 
        n192, sfr_wdat[5], n183, n176, n169, n163, n158}), .rdat({r_gpio_oe[1], 
        r_gpio_s1, r_gpio_oe[0], r_gpio_s0}) );
  glreg_8_00000032 u0_regD7 ( .clk(clk), .arstz(n79), .we(we_215), .wdat({n198, 
        n192, n188, n183, n177, n169, n165, n158}), .rdat({r_gpio_oe[3], 
        r_gpio_s3, r_gpio_oe[2], r_gpio_s2}) );
  glreg_a0_66 u0_regD9 ( .clk(clk), .arstz(n116), .we(we_217), .wdat({n198, 
        n192, sfr_wdat[5], n181, n177, n169, n163, n158}), .rdat({r_ana_tm, 
        r_fortxdat, r_fortxrdy, r_fortxen, r_sleep}) );
  glreg_a0_65 u0_regDE ( .clk(clk), .arstz(n115), .we(we_222), .wdat({n198, 
        n192, sfr_wdat[5], n181, n177, n169, n163, n158}), .rdat(regDE) );
  glsta_a0_3 u0_regDF ( .clk(clk), .arstz(n117), .rst0(1'b0), .set2(setDF), 
        .clr1(clrDF), .rdat(regDF), .irq(irqDF) );
  glreg_a0_64 u0_reg8F ( .clk(clk), .arstz(n113), .we(we_143), .wdat({n198, 
        n192, sfr_wdat[5], n181, n175, n169, n163, n158}), .rdat(r_dpdmctl) );
  glreg_WIDTH4 u0_reg94 ( .clk(clk), .arstz(n130), .we(we_148), .wdat({n192, 
        sfr_wdat[5], n181, n175}), .rdat(reg94[6:3]) );
  glreg_a0_63 u0_regA1 ( .clk(clk), .arstz(n111), .we(we[162]), .wdat({n198, 
        n192, sfr_wdat[5], n181, n175, n169, n163, n158}), .rdat(r_regtrm[7:0]) );
  glreg_a0_62 u0_regA2 ( .clk(clk), .arstz(n114), .we(we[162]), .wdat({n198, 
        n192, n188, n181, n175, n170, n163, n158}), .rdat(r_regtrm[15:8]) );
  glreg_a0_61 u0_regA3 ( .clk(clk), .arstz(n109), .we(we[163]), .wdat({n198, 
        n193, n188, n181, n175, n170, n163, n158}), .rdat(r_regtrm[23:16]) );
  glreg_a0_60 u0_regA4 ( .clk(clk), .arstz(n108), .we(we[164]), .wdat({n198, 
        n193, n187, n181, n175, n170, n164, n159}), .rdat(r_regtrm[31:24]) );
  glreg_a0_59 u0_regA5 ( .clk(clk), .arstz(n107), .we(we[165]), .wdat({n199, 
        n193, n187, n181, n175, n170, n164, n159}), .rdat(r_regtrm[39:32]) );
  glreg_a0_58 u0_regA6 ( .clk(clk), .arstz(n110), .we(we[166]), .wdat({n199, 
        n193, n187, n182, n175, n170, n164, n159}), .rdat(r_regtrm[47:40]) );
  glreg_a0_57 u0_regA7 ( .clk(clk), .arstz(n105), .we(we[167]), .wdat({n199, 
        n193, n187, n182, n175, n170, n164, n159}), .rdat(r_regtrm[55:48]) );
  glreg_a0_56 u0_regAB ( .clk(clk), .arstz(n104), .we(we_171), .wdat({n199, 
        n193, n187, n182, n175, n170, n164, n159}), .rdat(regAB) );
  glreg_8_00000028 u0_regAC ( .clk(clk), .arstz(n81), .we(we_172), .wdat({n199, 
        n193, n188, n182, n176, n170, n164, n159}), .rdat(regAC) );
  dbnc_WIDTH4_TIMEOUT14_2 u2_ovp_db ( .o_dbc(reg94[2]), .o_chg(), .i_org(
        srci[2]), .clk(clk_500), .rstz(n126) );
  dbnc_WIDTH4_TIMEOUT14_1 u1_ocp_db ( .o_dbc(reg94[1]), .o_chg(), .i_org(
        srci[1]), .clk(clk_500), .rstz(n125) );
  dbnc_WIDTH4_TIMEOUT14_0 u1_uvp_db ( .o_dbc(reg94[0]), .o_chg(), .i_org(
        srci[0]), .clk(clk_500), .rstz(n124) );
  dbnc_a0_2 u1_ovp_db ( .o_dbc(m_ovp), .o_chg(m_ovp_sta), .i_org(srci[2]), 
        .clk(clk_500k), .rstz(n123) );
  dbnc_WIDTH3_TIMEOUT5_4 u0_otpi_db ( .o_dbc(regAD[3]), .o_chg(setAE[3]), 
        .i_org(srci[5]), .clk(clk_1500k), .rstz(n128) );
  dbnc_WIDTH3_TIMEOUT5_3 u0_ocp_db ( .o_dbc(regAD[1]), .o_chg(setAE[1]), 
        .i_org(srci[1]), .clk(clk_1500k), .rstz(n129) );
  dbnc_WIDTH3_TIMEOUT5_2 u0_uvp_db ( .o_dbc(regAD[0]), .o_chg(setAE[0]), 
        .i_org(srci[0]), .clk(clk_1500k), .rstz(n127) );
  dbnc_WIDTH3_TIMEOUT5_1 u1_scp_db ( .o_dbc(m_scp), .o_chg(m_scp_sta), .i_org(
        srci[3]), .clk(clk_1500k), .rstz(n129) );
  dbnc_WIDTH3_TIMEOUT5_0 u0_dmf_db ( .o_dbc(regAD_7), .o_chg(setAE_7), .i_org(
        dm_fault), .clk(clk_1500k), .rstz(n128) );
  dbnc_WIDTH2_TIMEOUT2_13 u0_otps_db ( .o_dbc(reg94[7]), .o_chg(), .i_org(
        srci[5]), .clk(clk), .rstz(n131) );
  dbnc_WIDTH2_TIMEOUT2_12 u0_cc1_db ( .o_dbc(regF4_3), .o_chg(), .i_org(cc1_di), .clk(clk), .rstz(n131) );
  dbnc_WIDTH2_TIMEOUT2_11 u0_cc2_db ( .o_dbc(regF4_7_), .o_chg(), .i_org(
        cc2_di), .clk(clk), .rstz(n133) );
  dbnc_WIDTH2_TIMEOUT2_10 u0_ovp_db ( .o_dbc(s_ovp), .o_chg(s_ovp_sta), 
        .i_org(srci[2]), .clk(clk), .rstz(n133) );
  dbnc_WIDTH2_TIMEOUT2_9 u0_scp_db ( .o_dbc(s_scp), .o_chg(s_scp_sta), .i_org(
        srci[3]), .clk(clk), .rstz(n132) );
  dbnc_WIDTH2_TIMEOUT2_8 u0_v5oc_db ( .o_dbc(regAD[5]), .o_chg(setAE[5]), 
        .i_org(srci[4]), .clk(clk), .rstz(n132) );
  glsta_a0_2 u0_regAE ( .clk(clk), .arstz(n96), .rst0(1'b0), .set2({setAE_7, 
        1'b0, setAE}), .clr1(clrAE), .rdat(regAE), .irq(irqAE) );
  glreg_a0_55 u0_regAF ( .clk(clk), .arstz(n95), .we(we_175), .wdat({n199, 
        n193, n187, n182, n176, n170, n164, n159}), .rdat(regAF) );
  glreg_a0_54 u0_regE3 ( .clk(clk), .arstz(n102), .we(we_227), .wdat({n199, 
        n193, n187, n182, n176, n170, n164, n159}), .rdat({r_srcctl[7:4], 
        regE3, r_srcctl[1], regE3_0}) );
  glreg_4_00000004 u1_regE4 ( .clk(clk), .arstz(n130), .we(r_pwrv_upd), .wdat(
        lt_regE4_3_0), .rdat(r_fw_pwrv[3:0]) );
  glreg_8_00000004 u0_regE4 ( .clk(clk), .arstz(n84), .we(we_228), .wdat({n199, 
        n194, n187, n182, n176, n171, n164, n159}), .rdat({r_pwrctl, 
        lt_regE4_3_0}) );
  glreg_8_0000001f u0_regE5 ( .clk(clk), .arstz(n77), .we(r_pwrv_upd), .wdat({
        n199, n194, n188, n183, n177, n171, n165, n160}), .rdat(
        r_fw_pwrv[11:4]) );
  glreg_a0_53 u0_regE6 ( .clk(clk), .arstz(n98), .we(we_230), .wdat({n199, 
        n193, n187, n182, n176, n171, n164, n159}), .rdat(r_ccrx) );
  glreg_a0_52 u0_regE7 ( .clk(clk), .arstz(n91), .we(we_231), .wdat({n200, 
        n194, n188, n182, n176, n171, n165, n160}), .rdat(r_ccctl) );
  glreg_a0_51 u0_regE8 ( .clk(clk), .arstz(n90), .we(we_232), .wdat({n200, 
        n194, n188, n183, n176, n171, n165, n160}), .rdat(r_comp_opt) );
  glreg_a0_50 u0_regF5 ( .clk(clk), .arstz(n89), .we(we_245), .wdat({n200, 
        n194, n187, n182, n176, n171, n165, n160}), .rdat(r_cvctl) );
  glreg_a0_49 u0_regF6 ( .clk(clk), .arstz(n94), .we(we_246), .wdat({n198, 
        n192, n186, n180, n174, n168, sfr_wdat[1:0]}), .rdat(r_cctrx) );
  SNPS_CLOCK_GATE_HIGH_regbank_a0 clk_gate_rstcnt_reg ( .CLK(clk), .EN(N23), 
        .ENCLK(net10758), .TE(1'b0) );
  regbank_a0_DW01_add_0 add_527 ( .A(regAC), .B(regAB), .CI(1'b0), .SUM(
        r_pwr_i), .CO() );
  regbank_a0_DW01_inc_0 add_303 ( .A({1'b0, r_inst_ofs}), .SUM({
        SYNOPSYS_UNCONNECTED_1, inst_ofs_plus}) );
  regbank_a0_DW_rightsh_0 srl_132 ( .A({dac_r_vs, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, r_cctrx, r_cvctl, regF4_7_, x_daclsb[5:3], regF4_3, 
        x_daclsb[2:0], r_sar_en, r_dac_en, dac_r_ctl, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        r_comp_opt, r_ccctl, r_ccrx, r_fw_pwrv[11:4], r_pwrctl, r_fw_pwrv[3:0], 
        r_srcctl[7:4], regE3, r_srcctl[1], regE3_0, dac_r_cmpsta, dac_r_comp, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, regDF, regDE, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, r_ana_tm, r_fortxdat, 
        r_fortxrdy, r_fortxen, r_sleep, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, r_gpio_oe[3], r_gpio_s3, r_gpio_oe[2], r_gpio_s2, 
        r_gpio_oe[1], r_gpio_s1, r_gpio_oe[0], r_gpio_s0, r_gpio_pu[3:0], 
        r_gpio_pd[3:0], regD4, regD3_7_, r_gpio_oe[5], r_gpio_pu[5], 
        r_gpio_pd[5], regD3_3, r_gpio_oe[4], r_gpio_pu[4], r_gpio_pd[4], 
        i_i2c_rwbuf, r_exist1st, r_ordrs4, r_strtch, r_bclk_sel, r_gpio_tm, 
        r_gpio_oe[6], r_gpio_pu[6], r_gpio_pd[6], 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, reg31, reg30, i_i2c_ltbuf, reg28, reg27, r_i2c_deva, 
        r_hwi2c_en, 1'b0, 1'b0, r_i2c_attr, r_pg0_sel, reg25_0_, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, prx_rcvinf[4], REVID, 
        prx_rcvinf[3], ptx_fsm, prx_fsm, reg21, r_dat_portrole, r_dat_spec, 
        r_dat_datarole, reg20, reg19_7_, r_inst_ofs, i_i2c_ofs, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, dbgpo[31:24], r_auto_gdcrc[0], 
        r_auto_discard, r_spec, r_auto_gdcrc[1], prl_cpmsgid, prl_cany0, 
        prx_rcvinf[2:0], prl_fsm, reg12, r_txshrt, reg12_1, r_pshords, 
        reg11_7_, r_rxords_ena[6:5], reg11_4, r_rxords_ena[3:0], 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, pff_empty, 
        pff_full, pff_ptr, reg06, reg05, dbgpo[15:0], pff_rdat, r_last, 
        r_first, r_unlock, r_txnumk, r_txendk, r_txauto, regAF, regAE, regAD_7, 
        1'b0, regAD, regAC, regAB, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, r_regtrm, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, fcp_r_crc, fcp_r_dat, fcp_r_msk, fcp_r_sta, 
        fcp_r_ctl, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, fcp_r_acc, r_accctl, fcp_r_tui, reg94, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, r_isofs, r_adofs, r_dpdmctl, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, r_cvofs, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1}), .DATA_TC(1'b0), .SH({n155, sfr_addr[5:0], 
        1'b0, 1'b0, 1'b0}), .B({SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3, 
        SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6, 
        SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8, SYNOPSYS_UNCONNECTED_9, 
        SYNOPSYS_UNCONNECTED_10, SYNOPSYS_UNCONNECTED_11, 
        SYNOPSYS_UNCONNECTED_12, SYNOPSYS_UNCONNECTED_13, 
        SYNOPSYS_UNCONNECTED_14, SYNOPSYS_UNCONNECTED_15, 
        SYNOPSYS_UNCONNECTED_16, SYNOPSYS_UNCONNECTED_17, 
        SYNOPSYS_UNCONNECTED_18, SYNOPSYS_UNCONNECTED_19, 
        SYNOPSYS_UNCONNECTED_20, SYNOPSYS_UNCONNECTED_21, 
        SYNOPSYS_UNCONNECTED_22, SYNOPSYS_UNCONNECTED_23, 
        SYNOPSYS_UNCONNECTED_24, SYNOPSYS_UNCONNECTED_25, 
        SYNOPSYS_UNCONNECTED_26, SYNOPSYS_UNCONNECTED_27, 
        SYNOPSYS_UNCONNECTED_28, SYNOPSYS_UNCONNECTED_29, 
        SYNOPSYS_UNCONNECTED_30, SYNOPSYS_UNCONNECTED_31, 
        SYNOPSYS_UNCONNECTED_32, SYNOPSYS_UNCONNECTED_33, 
        SYNOPSYS_UNCONNECTED_34, SYNOPSYS_UNCONNECTED_35, 
        SYNOPSYS_UNCONNECTED_36, SYNOPSYS_UNCONNECTED_37, 
        SYNOPSYS_UNCONNECTED_38, SYNOPSYS_UNCONNECTED_39, 
        SYNOPSYS_UNCONNECTED_40, SYNOPSYS_UNCONNECTED_41, 
        SYNOPSYS_UNCONNECTED_42, SYNOPSYS_UNCONNECTED_43, 
        SYNOPSYS_UNCONNECTED_44, SYNOPSYS_UNCONNECTED_45, 
        SYNOPSYS_UNCONNECTED_46, SYNOPSYS_UNCONNECTED_47, 
        SYNOPSYS_UNCONNECTED_48, SYNOPSYS_UNCONNECTED_49, 
        SYNOPSYS_UNCONNECTED_50, SYNOPSYS_UNCONNECTED_51, 
        SYNOPSYS_UNCONNECTED_52, SYNOPSYS_UNCONNECTED_53, 
        SYNOPSYS_UNCONNECTED_54, SYNOPSYS_UNCONNECTED_55, 
        SYNOPSYS_UNCONNECTED_56, SYNOPSYS_UNCONNECTED_57, 
        SYNOPSYS_UNCONNECTED_58, SYNOPSYS_UNCONNECTED_59, 
        SYNOPSYS_UNCONNECTED_60, SYNOPSYS_UNCONNECTED_61, 
        SYNOPSYS_UNCONNECTED_62, SYNOPSYS_UNCONNECTED_63, 
        SYNOPSYS_UNCONNECTED_64, SYNOPSYS_UNCONNECTED_65, 
        SYNOPSYS_UNCONNECTED_66, SYNOPSYS_UNCONNECTED_67, 
        SYNOPSYS_UNCONNECTED_68, SYNOPSYS_UNCONNECTED_69, 
        SYNOPSYS_UNCONNECTED_70, SYNOPSYS_UNCONNECTED_71, 
        SYNOPSYS_UNCONNECTED_72, SYNOPSYS_UNCONNECTED_73, 
        SYNOPSYS_UNCONNECTED_74, SYNOPSYS_UNCONNECTED_75, 
        SYNOPSYS_UNCONNECTED_76, SYNOPSYS_UNCONNECTED_77, 
        SYNOPSYS_UNCONNECTED_78, SYNOPSYS_UNCONNECTED_79, 
        SYNOPSYS_UNCONNECTED_80, SYNOPSYS_UNCONNECTED_81, 
        SYNOPSYS_UNCONNECTED_82, SYNOPSYS_UNCONNECTED_83, 
        SYNOPSYS_UNCONNECTED_84, SYNOPSYS_UNCONNECTED_85, 
        SYNOPSYS_UNCONNECTED_86, SYNOPSYS_UNCONNECTED_87, 
        SYNOPSYS_UNCONNECTED_88, SYNOPSYS_UNCONNECTED_89, 
        SYNOPSYS_UNCONNECTED_90, SYNOPSYS_UNCONNECTED_91, 
        SYNOPSYS_UNCONNECTED_92, SYNOPSYS_UNCONNECTED_93, 
        SYNOPSYS_UNCONNECTED_94, SYNOPSYS_UNCONNECTED_95, 
        SYNOPSYS_UNCONNECTED_96, SYNOPSYS_UNCONNECTED_97, 
        SYNOPSYS_UNCONNECTED_98, SYNOPSYS_UNCONNECTED_99, 
        SYNOPSYS_UNCONNECTED_100, SYNOPSYS_UNCONNECTED_101, 
        SYNOPSYS_UNCONNECTED_102, SYNOPSYS_UNCONNECTED_103, 
        SYNOPSYS_UNCONNECTED_104, SYNOPSYS_UNCONNECTED_105, 
        SYNOPSYS_UNCONNECTED_106, SYNOPSYS_UNCONNECTED_107, 
        SYNOPSYS_UNCONNECTED_108, SYNOPSYS_UNCONNECTED_109, 
        SYNOPSYS_UNCONNECTED_110, SYNOPSYS_UNCONNECTED_111, 
        SYNOPSYS_UNCONNECTED_112, SYNOPSYS_UNCONNECTED_113, 
        SYNOPSYS_UNCONNECTED_114, SYNOPSYS_UNCONNECTED_115, 
        SYNOPSYS_UNCONNECTED_116, SYNOPSYS_UNCONNECTED_117, 
        SYNOPSYS_UNCONNECTED_118, SYNOPSYS_UNCONNECTED_119, 
        SYNOPSYS_UNCONNECTED_120, SYNOPSYS_UNCONNECTED_121, 
        SYNOPSYS_UNCONNECTED_122, SYNOPSYS_UNCONNECTED_123, 
        SYNOPSYS_UNCONNECTED_124, SYNOPSYS_UNCONNECTED_125, 
        SYNOPSYS_UNCONNECTED_126, SYNOPSYS_UNCONNECTED_127, 
        SYNOPSYS_UNCONNECTED_128, SYNOPSYS_UNCONNECTED_129, 
        SYNOPSYS_UNCONNECTED_130, SYNOPSYS_UNCONNECTED_131, 
        SYNOPSYS_UNCONNECTED_132, SYNOPSYS_UNCONNECTED_133, 
        SYNOPSYS_UNCONNECTED_134, SYNOPSYS_UNCONNECTED_135, 
        SYNOPSYS_UNCONNECTED_136, SYNOPSYS_UNCONNECTED_137, 
        SYNOPSYS_UNCONNECTED_138, SYNOPSYS_UNCONNECTED_139, 
        SYNOPSYS_UNCONNECTED_140, SYNOPSYS_UNCONNECTED_141, 
        SYNOPSYS_UNCONNECTED_142, SYNOPSYS_UNCONNECTED_143, 
        SYNOPSYS_UNCONNECTED_144, SYNOPSYS_UNCONNECTED_145, 
        SYNOPSYS_UNCONNECTED_146, SYNOPSYS_UNCONNECTED_147, 
        SYNOPSYS_UNCONNECTED_148, SYNOPSYS_UNCONNECTED_149, 
        SYNOPSYS_UNCONNECTED_150, SYNOPSYS_UNCONNECTED_151, 
        SYNOPSYS_UNCONNECTED_152, SYNOPSYS_UNCONNECTED_153, 
        SYNOPSYS_UNCONNECTED_154, SYNOPSYS_UNCONNECTED_155, 
        SYNOPSYS_UNCONNECTED_156, SYNOPSYS_UNCONNECTED_157, 
        SYNOPSYS_UNCONNECTED_158, SYNOPSYS_UNCONNECTED_159, 
        SYNOPSYS_UNCONNECTED_160, SYNOPSYS_UNCONNECTED_161, 
        SYNOPSYS_UNCONNECTED_162, SYNOPSYS_UNCONNECTED_163, 
        SYNOPSYS_UNCONNECTED_164, SYNOPSYS_UNCONNECTED_165, 
        SYNOPSYS_UNCONNECTED_166, SYNOPSYS_UNCONNECTED_167, 
        SYNOPSYS_UNCONNECTED_168, SYNOPSYS_UNCONNECTED_169, 
        SYNOPSYS_UNCONNECTED_170, SYNOPSYS_UNCONNECTED_171, 
        SYNOPSYS_UNCONNECTED_172, SYNOPSYS_UNCONNECTED_173, 
        SYNOPSYS_UNCONNECTED_174, SYNOPSYS_UNCONNECTED_175, 
        SYNOPSYS_UNCONNECTED_176, SYNOPSYS_UNCONNECTED_177, 
        SYNOPSYS_UNCONNECTED_178, SYNOPSYS_UNCONNECTED_179, 
        SYNOPSYS_UNCONNECTED_180, SYNOPSYS_UNCONNECTED_181, 
        SYNOPSYS_UNCONNECTED_182, SYNOPSYS_UNCONNECTED_183, 
        SYNOPSYS_UNCONNECTED_184, SYNOPSYS_UNCONNECTED_185, 
        SYNOPSYS_UNCONNECTED_186, SYNOPSYS_UNCONNECTED_187, 
        SYNOPSYS_UNCONNECTED_188, SYNOPSYS_UNCONNECTED_189, 
        SYNOPSYS_UNCONNECTED_190, SYNOPSYS_UNCONNECTED_191, 
        SYNOPSYS_UNCONNECTED_192, SYNOPSYS_UNCONNECTED_193, 
        SYNOPSYS_UNCONNECTED_194, SYNOPSYS_UNCONNECTED_195, 
        SYNOPSYS_UNCONNECTED_196, SYNOPSYS_UNCONNECTED_197, 
        SYNOPSYS_UNCONNECTED_198, SYNOPSYS_UNCONNECTED_199, 
        SYNOPSYS_UNCONNECTED_200, SYNOPSYS_UNCONNECTED_201, 
        SYNOPSYS_UNCONNECTED_202, SYNOPSYS_UNCONNECTED_203, 
        SYNOPSYS_UNCONNECTED_204, SYNOPSYS_UNCONNECTED_205, 
        SYNOPSYS_UNCONNECTED_206, SYNOPSYS_UNCONNECTED_207, 
        SYNOPSYS_UNCONNECTED_208, SYNOPSYS_UNCONNECTED_209, 
        SYNOPSYS_UNCONNECTED_210, SYNOPSYS_UNCONNECTED_211, 
        SYNOPSYS_UNCONNECTED_212, SYNOPSYS_UNCONNECTED_213, 
        SYNOPSYS_UNCONNECTED_214, SYNOPSYS_UNCONNECTED_215, 
        SYNOPSYS_UNCONNECTED_216, SYNOPSYS_UNCONNECTED_217, 
        SYNOPSYS_UNCONNECTED_218, SYNOPSYS_UNCONNECTED_219, 
        SYNOPSYS_UNCONNECTED_220, SYNOPSYS_UNCONNECTED_221, 
        SYNOPSYS_UNCONNECTED_222, SYNOPSYS_UNCONNECTED_223, 
        SYNOPSYS_UNCONNECTED_224, SYNOPSYS_UNCONNECTED_225, 
        SYNOPSYS_UNCONNECTED_226, SYNOPSYS_UNCONNECTED_227, 
        SYNOPSYS_UNCONNECTED_228, SYNOPSYS_UNCONNECTED_229, 
        SYNOPSYS_UNCONNECTED_230, SYNOPSYS_UNCONNECTED_231, 
        SYNOPSYS_UNCONNECTED_232, SYNOPSYS_UNCONNECTED_233, 
        SYNOPSYS_UNCONNECTED_234, SYNOPSYS_UNCONNECTED_235, 
        SYNOPSYS_UNCONNECTED_236, SYNOPSYS_UNCONNECTED_237, 
        SYNOPSYS_UNCONNECTED_238, SYNOPSYS_UNCONNECTED_239, 
        SYNOPSYS_UNCONNECTED_240, SYNOPSYS_UNCONNECTED_241, 
        SYNOPSYS_UNCONNECTED_242, SYNOPSYS_UNCONNECTED_243, 
        SYNOPSYS_UNCONNECTED_244, SYNOPSYS_UNCONNECTED_245, 
        SYNOPSYS_UNCONNECTED_246, SYNOPSYS_UNCONNECTED_247, 
        SYNOPSYS_UNCONNECTED_248, SYNOPSYS_UNCONNECTED_249, 
        SYNOPSYS_UNCONNECTED_250, SYNOPSYS_UNCONNECTED_251, 
        SYNOPSYS_UNCONNECTED_252, SYNOPSYS_UNCONNECTED_253, 
        SYNOPSYS_UNCONNECTED_254, SYNOPSYS_UNCONNECTED_255, 
        SYNOPSYS_UNCONNECTED_256, SYNOPSYS_UNCONNECTED_257, 
        SYNOPSYS_UNCONNECTED_258, SYNOPSYS_UNCONNECTED_259, 
        SYNOPSYS_UNCONNECTED_260, SYNOPSYS_UNCONNECTED_261, 
        SYNOPSYS_UNCONNECTED_262, SYNOPSYS_UNCONNECTED_263, 
        SYNOPSYS_UNCONNECTED_264, SYNOPSYS_UNCONNECTED_265, 
        SYNOPSYS_UNCONNECTED_266, SYNOPSYS_UNCONNECTED_267, 
        SYNOPSYS_UNCONNECTED_268, SYNOPSYS_UNCONNECTED_269, 
        SYNOPSYS_UNCONNECTED_270, SYNOPSYS_UNCONNECTED_271, 
        SYNOPSYS_UNCONNECTED_272, SYNOPSYS_UNCONNECTED_273, 
        SYNOPSYS_UNCONNECTED_274, SYNOPSYS_UNCONNECTED_275, 
        SYNOPSYS_UNCONNECTED_276, SYNOPSYS_UNCONNECTED_277, 
        SYNOPSYS_UNCONNECTED_278, SYNOPSYS_UNCONNECTED_279, 
        SYNOPSYS_UNCONNECTED_280, SYNOPSYS_UNCONNECTED_281, 
        SYNOPSYS_UNCONNECTED_282, SYNOPSYS_UNCONNECTED_283, 
        SYNOPSYS_UNCONNECTED_284, SYNOPSYS_UNCONNECTED_285, 
        SYNOPSYS_UNCONNECTED_286, SYNOPSYS_UNCONNECTED_287, 
        SYNOPSYS_UNCONNECTED_288, SYNOPSYS_UNCONNECTED_289, 
        SYNOPSYS_UNCONNECTED_290, SYNOPSYS_UNCONNECTED_291, 
        SYNOPSYS_UNCONNECTED_292, SYNOPSYS_UNCONNECTED_293, 
        SYNOPSYS_UNCONNECTED_294, SYNOPSYS_UNCONNECTED_295, 
        SYNOPSYS_UNCONNECTED_296, SYNOPSYS_UNCONNECTED_297, 
        SYNOPSYS_UNCONNECTED_298, SYNOPSYS_UNCONNECTED_299, 
        SYNOPSYS_UNCONNECTED_300, SYNOPSYS_UNCONNECTED_301, 
        SYNOPSYS_UNCONNECTED_302, SYNOPSYS_UNCONNECTED_303, 
        SYNOPSYS_UNCONNECTED_304, SYNOPSYS_UNCONNECTED_305, 
        SYNOPSYS_UNCONNECTED_306, SYNOPSYS_UNCONNECTED_307, 
        SYNOPSYS_UNCONNECTED_308, SYNOPSYS_UNCONNECTED_309, 
        SYNOPSYS_UNCONNECTED_310, SYNOPSYS_UNCONNECTED_311, 
        SYNOPSYS_UNCONNECTED_312, SYNOPSYS_UNCONNECTED_313, 
        SYNOPSYS_UNCONNECTED_314, SYNOPSYS_UNCONNECTED_315, 
        SYNOPSYS_UNCONNECTED_316, SYNOPSYS_UNCONNECTED_317, 
        SYNOPSYS_UNCONNECTED_318, SYNOPSYS_UNCONNECTED_319, 
        SYNOPSYS_UNCONNECTED_320, SYNOPSYS_UNCONNECTED_321, 
        SYNOPSYS_UNCONNECTED_322, SYNOPSYS_UNCONNECTED_323, 
        SYNOPSYS_UNCONNECTED_324, SYNOPSYS_UNCONNECTED_325, 
        SYNOPSYS_UNCONNECTED_326, SYNOPSYS_UNCONNECTED_327, 
        SYNOPSYS_UNCONNECTED_328, SYNOPSYS_UNCONNECTED_329, 
        SYNOPSYS_UNCONNECTED_330, SYNOPSYS_UNCONNECTED_331, 
        SYNOPSYS_UNCONNECTED_332, SYNOPSYS_UNCONNECTED_333, 
        SYNOPSYS_UNCONNECTED_334, SYNOPSYS_UNCONNECTED_335, 
        SYNOPSYS_UNCONNECTED_336, SYNOPSYS_UNCONNECTED_337, 
        SYNOPSYS_UNCONNECTED_338, SYNOPSYS_UNCONNECTED_339, 
        SYNOPSYS_UNCONNECTED_340, SYNOPSYS_UNCONNECTED_341, 
        SYNOPSYS_UNCONNECTED_342, SYNOPSYS_UNCONNECTED_343, 
        SYNOPSYS_UNCONNECTED_344, SYNOPSYS_UNCONNECTED_345, 
        SYNOPSYS_UNCONNECTED_346, SYNOPSYS_UNCONNECTED_347, 
        SYNOPSYS_UNCONNECTED_348, SYNOPSYS_UNCONNECTED_349, 
        SYNOPSYS_UNCONNECTED_350, SYNOPSYS_UNCONNECTED_351, 
        SYNOPSYS_UNCONNECTED_352, SYNOPSYS_UNCONNECTED_353, 
        SYNOPSYS_UNCONNECTED_354, SYNOPSYS_UNCONNECTED_355, 
        SYNOPSYS_UNCONNECTED_356, SYNOPSYS_UNCONNECTED_357, 
        SYNOPSYS_UNCONNECTED_358, SYNOPSYS_UNCONNECTED_359, 
        SYNOPSYS_UNCONNECTED_360, SYNOPSYS_UNCONNECTED_361, 
        SYNOPSYS_UNCONNECTED_362, SYNOPSYS_UNCONNECTED_363, 
        SYNOPSYS_UNCONNECTED_364, SYNOPSYS_UNCONNECTED_365, 
        SYNOPSYS_UNCONNECTED_366, SYNOPSYS_UNCONNECTED_367, 
        SYNOPSYS_UNCONNECTED_368, SYNOPSYS_UNCONNECTED_369, 
        SYNOPSYS_UNCONNECTED_370, SYNOPSYS_UNCONNECTED_371, 
        SYNOPSYS_UNCONNECTED_372, SYNOPSYS_UNCONNECTED_373, 
        SYNOPSYS_UNCONNECTED_374, SYNOPSYS_UNCONNECTED_375, 
        SYNOPSYS_UNCONNECTED_376, SYNOPSYS_UNCONNECTED_377, 
        SYNOPSYS_UNCONNECTED_378, SYNOPSYS_UNCONNECTED_379, 
        SYNOPSYS_UNCONNECTED_380, SYNOPSYS_UNCONNECTED_381, 
        SYNOPSYS_UNCONNECTED_382, SYNOPSYS_UNCONNECTED_383, 
        SYNOPSYS_UNCONNECTED_384, SYNOPSYS_UNCONNECTED_385, 
        SYNOPSYS_UNCONNECTED_386, SYNOPSYS_UNCONNECTED_387, 
        SYNOPSYS_UNCONNECTED_388, SYNOPSYS_UNCONNECTED_389, 
        SYNOPSYS_UNCONNECTED_390, SYNOPSYS_UNCONNECTED_391, 
        SYNOPSYS_UNCONNECTED_392, SYNOPSYS_UNCONNECTED_393, 
        SYNOPSYS_UNCONNECTED_394, SYNOPSYS_UNCONNECTED_395, 
        SYNOPSYS_UNCONNECTED_396, SYNOPSYS_UNCONNECTED_397, 
        SYNOPSYS_UNCONNECTED_398, SYNOPSYS_UNCONNECTED_399, 
        SYNOPSYS_UNCONNECTED_400, SYNOPSYS_UNCONNECTED_401, 
        SYNOPSYS_UNCONNECTED_402, SYNOPSYS_UNCONNECTED_403, 
        SYNOPSYS_UNCONNECTED_404, SYNOPSYS_UNCONNECTED_405, 
        SYNOPSYS_UNCONNECTED_406, SYNOPSYS_UNCONNECTED_407, 
        SYNOPSYS_UNCONNECTED_408, SYNOPSYS_UNCONNECTED_409, 
        SYNOPSYS_UNCONNECTED_410, SYNOPSYS_UNCONNECTED_411, 
        SYNOPSYS_UNCONNECTED_412, SYNOPSYS_UNCONNECTED_413, 
        SYNOPSYS_UNCONNECTED_414, SYNOPSYS_UNCONNECTED_415, 
        SYNOPSYS_UNCONNECTED_416, SYNOPSYS_UNCONNECTED_417, 
        SYNOPSYS_UNCONNECTED_418, SYNOPSYS_UNCONNECTED_419, 
        SYNOPSYS_UNCONNECTED_420, SYNOPSYS_UNCONNECTED_421, 
        SYNOPSYS_UNCONNECTED_422, SYNOPSYS_UNCONNECTED_423, 
        SYNOPSYS_UNCONNECTED_424, SYNOPSYS_UNCONNECTED_425, 
        SYNOPSYS_UNCONNECTED_426, SYNOPSYS_UNCONNECTED_427, 
        SYNOPSYS_UNCONNECTED_428, SYNOPSYS_UNCONNECTED_429, 
        SYNOPSYS_UNCONNECTED_430, SYNOPSYS_UNCONNECTED_431, 
        SYNOPSYS_UNCONNECTED_432, SYNOPSYS_UNCONNECTED_433, 
        SYNOPSYS_UNCONNECTED_434, SYNOPSYS_UNCONNECTED_435, 
        SYNOPSYS_UNCONNECTED_436, SYNOPSYS_UNCONNECTED_437, 
        SYNOPSYS_UNCONNECTED_438, SYNOPSYS_UNCONNECTED_439, 
        SYNOPSYS_UNCONNECTED_440, SYNOPSYS_UNCONNECTED_441, 
        SYNOPSYS_UNCONNECTED_442, SYNOPSYS_UNCONNECTED_443, 
        SYNOPSYS_UNCONNECTED_444, SYNOPSYS_UNCONNECTED_445, 
        SYNOPSYS_UNCONNECTED_446, SYNOPSYS_UNCONNECTED_447, 
        SYNOPSYS_UNCONNECTED_448, SYNOPSYS_UNCONNECTED_449, 
        SYNOPSYS_UNCONNECTED_450, SYNOPSYS_UNCONNECTED_451, 
        SYNOPSYS_UNCONNECTED_452, SYNOPSYS_UNCONNECTED_453, 
        SYNOPSYS_UNCONNECTED_454, SYNOPSYS_UNCONNECTED_455, 
        SYNOPSYS_UNCONNECTED_456, SYNOPSYS_UNCONNECTED_457, 
        SYNOPSYS_UNCONNECTED_458, SYNOPSYS_UNCONNECTED_459, 
        SYNOPSYS_UNCONNECTED_460, SYNOPSYS_UNCONNECTED_461, 
        SYNOPSYS_UNCONNECTED_462, SYNOPSYS_UNCONNECTED_463, 
        SYNOPSYS_UNCONNECTED_464, SYNOPSYS_UNCONNECTED_465, 
        SYNOPSYS_UNCONNECTED_466, SYNOPSYS_UNCONNECTED_467, 
        SYNOPSYS_UNCONNECTED_468, SYNOPSYS_UNCONNECTED_469, 
        SYNOPSYS_UNCONNECTED_470, SYNOPSYS_UNCONNECTED_471, 
        SYNOPSYS_UNCONNECTED_472, SYNOPSYS_UNCONNECTED_473, 
        SYNOPSYS_UNCONNECTED_474, SYNOPSYS_UNCONNECTED_475, 
        SYNOPSYS_UNCONNECTED_476, SYNOPSYS_UNCONNECTED_477, 
        SYNOPSYS_UNCONNECTED_478, SYNOPSYS_UNCONNECTED_479, 
        SYNOPSYS_UNCONNECTED_480, SYNOPSYS_UNCONNECTED_481, 
        SYNOPSYS_UNCONNECTED_482, SYNOPSYS_UNCONNECTED_483, 
        SYNOPSYS_UNCONNECTED_484, SYNOPSYS_UNCONNECTED_485, 
        SYNOPSYS_UNCONNECTED_486, SYNOPSYS_UNCONNECTED_487, 
        SYNOPSYS_UNCONNECTED_488, SYNOPSYS_UNCONNECTED_489, 
        SYNOPSYS_UNCONNECTED_490, SYNOPSYS_UNCONNECTED_491, 
        SYNOPSYS_UNCONNECTED_492, SYNOPSYS_UNCONNECTED_493, 
        SYNOPSYS_UNCONNECTED_494, SYNOPSYS_UNCONNECTED_495, 
        SYNOPSYS_UNCONNECTED_496, SYNOPSYS_UNCONNECTED_497, 
        SYNOPSYS_UNCONNECTED_498, SYNOPSYS_UNCONNECTED_499, 
        SYNOPSYS_UNCONNECTED_500, SYNOPSYS_UNCONNECTED_501, 
        SYNOPSYS_UNCONNECTED_502, SYNOPSYS_UNCONNECTED_503, 
        SYNOPSYS_UNCONNECTED_504, SYNOPSYS_UNCONNECTED_505, 
        SYNOPSYS_UNCONNECTED_506, SYNOPSYS_UNCONNECTED_507, 
        SYNOPSYS_UNCONNECTED_508, SYNOPSYS_UNCONNECTED_509, 
        SYNOPSYS_UNCONNECTED_510, SYNOPSYS_UNCONNECTED_511, 
        SYNOPSYS_UNCONNECTED_512, SYNOPSYS_UNCONNECTED_513, 
        SYNOPSYS_UNCONNECTED_514, SYNOPSYS_UNCONNECTED_515, 
        SYNOPSYS_UNCONNECTED_516, SYNOPSYS_UNCONNECTED_517, 
        SYNOPSYS_UNCONNECTED_518, SYNOPSYS_UNCONNECTED_519, 
        SYNOPSYS_UNCONNECTED_520, SYNOPSYS_UNCONNECTED_521, 
        SYNOPSYS_UNCONNECTED_522, SYNOPSYS_UNCONNECTED_523, 
        SYNOPSYS_UNCONNECTED_524, SYNOPSYS_UNCONNECTED_525, 
        SYNOPSYS_UNCONNECTED_526, SYNOPSYS_UNCONNECTED_527, 
        SYNOPSYS_UNCONNECTED_528, SYNOPSYS_UNCONNECTED_529, 
        SYNOPSYS_UNCONNECTED_530, SYNOPSYS_UNCONNECTED_531, 
        SYNOPSYS_UNCONNECTED_532, SYNOPSYS_UNCONNECTED_533, 
        SYNOPSYS_UNCONNECTED_534, SYNOPSYS_UNCONNECTED_535, 
        SYNOPSYS_UNCONNECTED_536, SYNOPSYS_UNCONNECTED_537, 
        SYNOPSYS_UNCONNECTED_538, SYNOPSYS_UNCONNECTED_539, 
        SYNOPSYS_UNCONNECTED_540, SYNOPSYS_UNCONNECTED_541, 
        SYNOPSYS_UNCONNECTED_542, SYNOPSYS_UNCONNECTED_543, 
        SYNOPSYS_UNCONNECTED_544, SYNOPSYS_UNCONNECTED_545, 
        SYNOPSYS_UNCONNECTED_546, SYNOPSYS_UNCONNECTED_547, 
        SYNOPSYS_UNCONNECTED_548, SYNOPSYS_UNCONNECTED_549, 
        SYNOPSYS_UNCONNECTED_550, SYNOPSYS_UNCONNECTED_551, 
        SYNOPSYS_UNCONNECTED_552, SYNOPSYS_UNCONNECTED_553, 
        SYNOPSYS_UNCONNECTED_554, SYNOPSYS_UNCONNECTED_555, 
        SYNOPSYS_UNCONNECTED_556, SYNOPSYS_UNCONNECTED_557, 
        SYNOPSYS_UNCONNECTED_558, SYNOPSYS_UNCONNECTED_559, 
        SYNOPSYS_UNCONNECTED_560, SYNOPSYS_UNCONNECTED_561, 
        SYNOPSYS_UNCONNECTED_562, SYNOPSYS_UNCONNECTED_563, 
        SYNOPSYS_UNCONNECTED_564, SYNOPSYS_UNCONNECTED_565, 
        SYNOPSYS_UNCONNECTED_566, SYNOPSYS_UNCONNECTED_567, 
        SYNOPSYS_UNCONNECTED_568, SYNOPSYS_UNCONNECTED_569, 
        SYNOPSYS_UNCONNECTED_570, SYNOPSYS_UNCONNECTED_571, 
        SYNOPSYS_UNCONNECTED_572, SYNOPSYS_UNCONNECTED_573, 
        SYNOPSYS_UNCONNECTED_574, SYNOPSYS_UNCONNECTED_575, 
        SYNOPSYS_UNCONNECTED_576, SYNOPSYS_UNCONNECTED_577, 
        SYNOPSYS_UNCONNECTED_578, SYNOPSYS_UNCONNECTED_579, 
        SYNOPSYS_UNCONNECTED_580, SYNOPSYS_UNCONNECTED_581, 
        SYNOPSYS_UNCONNECTED_582, SYNOPSYS_UNCONNECTED_583, 
        SYNOPSYS_UNCONNECTED_584, SYNOPSYS_UNCONNECTED_585, 
        SYNOPSYS_UNCONNECTED_586, SYNOPSYS_UNCONNECTED_587, 
        SYNOPSYS_UNCONNECTED_588, SYNOPSYS_UNCONNECTED_589, 
        SYNOPSYS_UNCONNECTED_590, SYNOPSYS_UNCONNECTED_591, 
        SYNOPSYS_UNCONNECTED_592, SYNOPSYS_UNCONNECTED_593, 
        SYNOPSYS_UNCONNECTED_594, SYNOPSYS_UNCONNECTED_595, 
        SYNOPSYS_UNCONNECTED_596, SYNOPSYS_UNCONNECTED_597, 
        SYNOPSYS_UNCONNECTED_598, SYNOPSYS_UNCONNECTED_599, 
        SYNOPSYS_UNCONNECTED_600, SYNOPSYS_UNCONNECTED_601, 
        SYNOPSYS_UNCONNECTED_602, SYNOPSYS_UNCONNECTED_603, 
        SYNOPSYS_UNCONNECTED_604, SYNOPSYS_UNCONNECTED_605, 
        SYNOPSYS_UNCONNECTED_606, SYNOPSYS_UNCONNECTED_607, 
        SYNOPSYS_UNCONNECTED_608, SYNOPSYS_UNCONNECTED_609, 
        SYNOPSYS_UNCONNECTED_610, SYNOPSYS_UNCONNECTED_611, 
        SYNOPSYS_UNCONNECTED_612, SYNOPSYS_UNCONNECTED_613, 
        SYNOPSYS_UNCONNECTED_614, SYNOPSYS_UNCONNECTED_615, 
        SYNOPSYS_UNCONNECTED_616, SYNOPSYS_UNCONNECTED_617, 
        SYNOPSYS_UNCONNECTED_618, SYNOPSYS_UNCONNECTED_619, 
        SYNOPSYS_UNCONNECTED_620, SYNOPSYS_UNCONNECTED_621, 
        SYNOPSYS_UNCONNECTED_622, SYNOPSYS_UNCONNECTED_623, 
        SYNOPSYS_UNCONNECTED_624, SYNOPSYS_UNCONNECTED_625, 
        SYNOPSYS_UNCONNECTED_626, SYNOPSYS_UNCONNECTED_627, 
        SYNOPSYS_UNCONNECTED_628, SYNOPSYS_UNCONNECTED_629, 
        SYNOPSYS_UNCONNECTED_630, SYNOPSYS_UNCONNECTED_631, 
        SYNOPSYS_UNCONNECTED_632, SYNOPSYS_UNCONNECTED_633, 
        SYNOPSYS_UNCONNECTED_634, SYNOPSYS_UNCONNECTED_635, 
        SYNOPSYS_UNCONNECTED_636, SYNOPSYS_UNCONNECTED_637, 
        SYNOPSYS_UNCONNECTED_638, SYNOPSYS_UNCONNECTED_639, 
        SYNOPSYS_UNCONNECTED_640, SYNOPSYS_UNCONNECTED_641, 
        SYNOPSYS_UNCONNECTED_642, SYNOPSYS_UNCONNECTED_643, 
        SYNOPSYS_UNCONNECTED_644, SYNOPSYS_UNCONNECTED_645, 
        SYNOPSYS_UNCONNECTED_646, SYNOPSYS_UNCONNECTED_647, 
        SYNOPSYS_UNCONNECTED_648, SYNOPSYS_UNCONNECTED_649, 
        SYNOPSYS_UNCONNECTED_650, SYNOPSYS_UNCONNECTED_651, 
        SYNOPSYS_UNCONNECTED_652, SYNOPSYS_UNCONNECTED_653, 
        SYNOPSYS_UNCONNECTED_654, SYNOPSYS_UNCONNECTED_655, 
        SYNOPSYS_UNCONNECTED_656, SYNOPSYS_UNCONNECTED_657, 
        SYNOPSYS_UNCONNECTED_658, SYNOPSYS_UNCONNECTED_659, 
        SYNOPSYS_UNCONNECTED_660, SYNOPSYS_UNCONNECTED_661, 
        SYNOPSYS_UNCONNECTED_662, SYNOPSYS_UNCONNECTED_663, 
        SYNOPSYS_UNCONNECTED_664, SYNOPSYS_UNCONNECTED_665, 
        SYNOPSYS_UNCONNECTED_666, SYNOPSYS_UNCONNECTED_667, 
        SYNOPSYS_UNCONNECTED_668, SYNOPSYS_UNCONNECTED_669, 
        SYNOPSYS_UNCONNECTED_670, SYNOPSYS_UNCONNECTED_671, 
        SYNOPSYS_UNCONNECTED_672, SYNOPSYS_UNCONNECTED_673, 
        SYNOPSYS_UNCONNECTED_674, SYNOPSYS_UNCONNECTED_675, 
        SYNOPSYS_UNCONNECTED_676, SYNOPSYS_UNCONNECTED_677, 
        SYNOPSYS_UNCONNECTED_678, SYNOPSYS_UNCONNECTED_679, 
        SYNOPSYS_UNCONNECTED_680, SYNOPSYS_UNCONNECTED_681, 
        SYNOPSYS_UNCONNECTED_682, SYNOPSYS_UNCONNECTED_683, 
        SYNOPSYS_UNCONNECTED_684, SYNOPSYS_UNCONNECTED_685, 
        SYNOPSYS_UNCONNECTED_686, SYNOPSYS_UNCONNECTED_687, 
        SYNOPSYS_UNCONNECTED_688, SYNOPSYS_UNCONNECTED_689, 
        SYNOPSYS_UNCONNECTED_690, SYNOPSYS_UNCONNECTED_691, 
        SYNOPSYS_UNCONNECTED_692, SYNOPSYS_UNCONNECTED_693, 
        SYNOPSYS_UNCONNECTED_694, SYNOPSYS_UNCONNECTED_695, 
        SYNOPSYS_UNCONNECTED_696, SYNOPSYS_UNCONNECTED_697, 
        SYNOPSYS_UNCONNECTED_698, SYNOPSYS_UNCONNECTED_699, 
        SYNOPSYS_UNCONNECTED_700, SYNOPSYS_UNCONNECTED_701, 
        SYNOPSYS_UNCONNECTED_702, SYNOPSYS_UNCONNECTED_703, 
        SYNOPSYS_UNCONNECTED_704, SYNOPSYS_UNCONNECTED_705, 
        SYNOPSYS_UNCONNECTED_706, SYNOPSYS_UNCONNECTED_707, 
        SYNOPSYS_UNCONNECTED_708, SYNOPSYS_UNCONNECTED_709, 
        SYNOPSYS_UNCONNECTED_710, SYNOPSYS_UNCONNECTED_711, 
        SYNOPSYS_UNCONNECTED_712, SYNOPSYS_UNCONNECTED_713, 
        SYNOPSYS_UNCONNECTED_714, SYNOPSYS_UNCONNECTED_715, 
        SYNOPSYS_UNCONNECTED_716, SYNOPSYS_UNCONNECTED_717, 
        SYNOPSYS_UNCONNECTED_718, SYNOPSYS_UNCONNECTED_719, 
        SYNOPSYS_UNCONNECTED_720, SYNOPSYS_UNCONNECTED_721, 
        SYNOPSYS_UNCONNECTED_722, SYNOPSYS_UNCONNECTED_723, 
        SYNOPSYS_UNCONNECTED_724, SYNOPSYS_UNCONNECTED_725, 
        SYNOPSYS_UNCONNECTED_726, SYNOPSYS_UNCONNECTED_727, 
        SYNOPSYS_UNCONNECTED_728, SYNOPSYS_UNCONNECTED_729, 
        SYNOPSYS_UNCONNECTED_730, SYNOPSYS_UNCONNECTED_731, 
        SYNOPSYS_UNCONNECTED_732, SYNOPSYS_UNCONNECTED_733, 
        SYNOPSYS_UNCONNECTED_734, SYNOPSYS_UNCONNECTED_735, 
        SYNOPSYS_UNCONNECTED_736, SYNOPSYS_UNCONNECTED_737, 
        SYNOPSYS_UNCONNECTED_738, SYNOPSYS_UNCONNECTED_739, 
        SYNOPSYS_UNCONNECTED_740, SYNOPSYS_UNCONNECTED_741, 
        SYNOPSYS_UNCONNECTED_742, SYNOPSYS_UNCONNECTED_743, 
        SYNOPSYS_UNCONNECTED_744, SYNOPSYS_UNCONNECTED_745, 
        SYNOPSYS_UNCONNECTED_746, SYNOPSYS_UNCONNECTED_747, 
        SYNOPSYS_UNCONNECTED_748, SYNOPSYS_UNCONNECTED_749, 
        SYNOPSYS_UNCONNECTED_750, SYNOPSYS_UNCONNECTED_751, 
        SYNOPSYS_UNCONNECTED_752, SYNOPSYS_UNCONNECTED_753, 
        SYNOPSYS_UNCONNECTED_754, SYNOPSYS_UNCONNECTED_755, 
        SYNOPSYS_UNCONNECTED_756, SYNOPSYS_UNCONNECTED_757, 
        SYNOPSYS_UNCONNECTED_758, SYNOPSYS_UNCONNECTED_759, 
        SYNOPSYS_UNCONNECTED_760, SYNOPSYS_UNCONNECTED_761, 
        SYNOPSYS_UNCONNECTED_762, SYNOPSYS_UNCONNECTED_763, 
        SYNOPSYS_UNCONNECTED_764, SYNOPSYS_UNCONNECTED_765, 
        SYNOPSYS_UNCONNECTED_766, SYNOPSYS_UNCONNECTED_767, 
        SYNOPSYS_UNCONNECTED_768, SYNOPSYS_UNCONNECTED_769, 
        SYNOPSYS_UNCONNECTED_770, SYNOPSYS_UNCONNECTED_771, 
        SYNOPSYS_UNCONNECTED_772, SYNOPSYS_UNCONNECTED_773, 
        SYNOPSYS_UNCONNECTED_774, SYNOPSYS_UNCONNECTED_775, 
        SYNOPSYS_UNCONNECTED_776, SYNOPSYS_UNCONNECTED_777, 
        SYNOPSYS_UNCONNECTED_778, SYNOPSYS_UNCONNECTED_779, 
        SYNOPSYS_UNCONNECTED_780, SYNOPSYS_UNCONNECTED_781, 
        SYNOPSYS_UNCONNECTED_782, SYNOPSYS_UNCONNECTED_783, 
        SYNOPSYS_UNCONNECTED_784, SYNOPSYS_UNCONNECTED_785, 
        SYNOPSYS_UNCONNECTED_786, SYNOPSYS_UNCONNECTED_787, 
        SYNOPSYS_UNCONNECTED_788, SYNOPSYS_UNCONNECTED_789, 
        SYNOPSYS_UNCONNECTED_790, SYNOPSYS_UNCONNECTED_791, 
        SYNOPSYS_UNCONNECTED_792, SYNOPSYS_UNCONNECTED_793, 
        SYNOPSYS_UNCONNECTED_794, SYNOPSYS_UNCONNECTED_795, 
        SYNOPSYS_UNCONNECTED_796, SYNOPSYS_UNCONNECTED_797, 
        SYNOPSYS_UNCONNECTED_798, SYNOPSYS_UNCONNECTED_799, 
        SYNOPSYS_UNCONNECTED_800, SYNOPSYS_UNCONNECTED_801, 
        SYNOPSYS_UNCONNECTED_802, SYNOPSYS_UNCONNECTED_803, 
        SYNOPSYS_UNCONNECTED_804, SYNOPSYS_UNCONNECTED_805, 
        SYNOPSYS_UNCONNECTED_806, SYNOPSYS_UNCONNECTED_807, 
        SYNOPSYS_UNCONNECTED_808, SYNOPSYS_UNCONNECTED_809, 
        SYNOPSYS_UNCONNECTED_810, SYNOPSYS_UNCONNECTED_811, 
        SYNOPSYS_UNCONNECTED_812, SYNOPSYS_UNCONNECTED_813, 
        SYNOPSYS_UNCONNECTED_814, SYNOPSYS_UNCONNECTED_815, 
        SYNOPSYS_UNCONNECTED_816, SYNOPSYS_UNCONNECTED_817, 
        SYNOPSYS_UNCONNECTED_818, SYNOPSYS_UNCONNECTED_819, 
        SYNOPSYS_UNCONNECTED_820, SYNOPSYS_UNCONNECTED_821, 
        SYNOPSYS_UNCONNECTED_822, SYNOPSYS_UNCONNECTED_823, 
        SYNOPSYS_UNCONNECTED_824, SYNOPSYS_UNCONNECTED_825, 
        SYNOPSYS_UNCONNECTED_826, SYNOPSYS_UNCONNECTED_827, 
        SYNOPSYS_UNCONNECTED_828, SYNOPSYS_UNCONNECTED_829, 
        SYNOPSYS_UNCONNECTED_830, SYNOPSYS_UNCONNECTED_831, 
        SYNOPSYS_UNCONNECTED_832, SYNOPSYS_UNCONNECTED_833, 
        SYNOPSYS_UNCONNECTED_834, SYNOPSYS_UNCONNECTED_835, 
        SYNOPSYS_UNCONNECTED_836, SYNOPSYS_UNCONNECTED_837, 
        SYNOPSYS_UNCONNECTED_838, SYNOPSYS_UNCONNECTED_839, 
        SYNOPSYS_UNCONNECTED_840, SYNOPSYS_UNCONNECTED_841, 
        SYNOPSYS_UNCONNECTED_842, SYNOPSYS_UNCONNECTED_843, 
        SYNOPSYS_UNCONNECTED_844, SYNOPSYS_UNCONNECTED_845, 
        SYNOPSYS_UNCONNECTED_846, SYNOPSYS_UNCONNECTED_847, 
        SYNOPSYS_UNCONNECTED_848, SYNOPSYS_UNCONNECTED_849, 
        SYNOPSYS_UNCONNECTED_850, SYNOPSYS_UNCONNECTED_851, 
        SYNOPSYS_UNCONNECTED_852, SYNOPSYS_UNCONNECTED_853, 
        SYNOPSYS_UNCONNECTED_854, SYNOPSYS_UNCONNECTED_855, 
        SYNOPSYS_UNCONNECTED_856, SYNOPSYS_UNCONNECTED_857, 
        SYNOPSYS_UNCONNECTED_858, SYNOPSYS_UNCONNECTED_859, 
        SYNOPSYS_UNCONNECTED_860, SYNOPSYS_UNCONNECTED_861, 
        SYNOPSYS_UNCONNECTED_862, SYNOPSYS_UNCONNECTED_863, 
        SYNOPSYS_UNCONNECTED_864, SYNOPSYS_UNCONNECTED_865, 
        SYNOPSYS_UNCONNECTED_866, SYNOPSYS_UNCONNECTED_867, 
        SYNOPSYS_UNCONNECTED_868, SYNOPSYS_UNCONNECTED_869, 
        SYNOPSYS_UNCONNECTED_870, SYNOPSYS_UNCONNECTED_871, 
        SYNOPSYS_UNCONNECTED_872, SYNOPSYS_UNCONNECTED_873, 
        SYNOPSYS_UNCONNECTED_874, SYNOPSYS_UNCONNECTED_875, 
        SYNOPSYS_UNCONNECTED_876, SYNOPSYS_UNCONNECTED_877, 
        SYNOPSYS_UNCONNECTED_878, SYNOPSYS_UNCONNECTED_879, 
        SYNOPSYS_UNCONNECTED_880, SYNOPSYS_UNCONNECTED_881, 
        SYNOPSYS_UNCONNECTED_882, SYNOPSYS_UNCONNECTED_883, 
        SYNOPSYS_UNCONNECTED_884, SYNOPSYS_UNCONNECTED_885, 
        SYNOPSYS_UNCONNECTED_886, SYNOPSYS_UNCONNECTED_887, 
        SYNOPSYS_UNCONNECTED_888, SYNOPSYS_UNCONNECTED_889, 
        SYNOPSYS_UNCONNECTED_890, SYNOPSYS_UNCONNECTED_891, 
        SYNOPSYS_UNCONNECTED_892, SYNOPSYS_UNCONNECTED_893, 
        SYNOPSYS_UNCONNECTED_894, SYNOPSYS_UNCONNECTED_895, 
        SYNOPSYS_UNCONNECTED_896, SYNOPSYS_UNCONNECTED_897, 
        SYNOPSYS_UNCONNECTED_898, SYNOPSYS_UNCONNECTED_899, 
        SYNOPSYS_UNCONNECTED_900, SYNOPSYS_UNCONNECTED_901, 
        SYNOPSYS_UNCONNECTED_902, SYNOPSYS_UNCONNECTED_903, 
        SYNOPSYS_UNCONNECTED_904, SYNOPSYS_UNCONNECTED_905, 
        SYNOPSYS_UNCONNECTED_906, SYNOPSYS_UNCONNECTED_907, 
        SYNOPSYS_UNCONNECTED_908, SYNOPSYS_UNCONNECTED_909, 
        SYNOPSYS_UNCONNECTED_910, SYNOPSYS_UNCONNECTED_911, 
        SYNOPSYS_UNCONNECTED_912, SYNOPSYS_UNCONNECTED_913, 
        SYNOPSYS_UNCONNECTED_914, SYNOPSYS_UNCONNECTED_915, 
        SYNOPSYS_UNCONNECTED_916, SYNOPSYS_UNCONNECTED_917, 
        SYNOPSYS_UNCONNECTED_918, SYNOPSYS_UNCONNECTED_919, 
        SYNOPSYS_UNCONNECTED_920, SYNOPSYS_UNCONNECTED_921, 
        SYNOPSYS_UNCONNECTED_922, SYNOPSYS_UNCONNECTED_923, 
        SYNOPSYS_UNCONNECTED_924, SYNOPSYS_UNCONNECTED_925, 
        SYNOPSYS_UNCONNECTED_926, SYNOPSYS_UNCONNECTED_927, 
        SYNOPSYS_UNCONNECTED_928, SYNOPSYS_UNCONNECTED_929, 
        SYNOPSYS_UNCONNECTED_930, SYNOPSYS_UNCONNECTED_931, 
        SYNOPSYS_UNCONNECTED_932, SYNOPSYS_UNCONNECTED_933, 
        SYNOPSYS_UNCONNECTED_934, SYNOPSYS_UNCONNECTED_935, 
        SYNOPSYS_UNCONNECTED_936, SYNOPSYS_UNCONNECTED_937, 
        SYNOPSYS_UNCONNECTED_938, SYNOPSYS_UNCONNECTED_939, 
        SYNOPSYS_UNCONNECTED_940, SYNOPSYS_UNCONNECTED_941, 
        SYNOPSYS_UNCONNECTED_942, SYNOPSYS_UNCONNECTED_943, 
        SYNOPSYS_UNCONNECTED_944, SYNOPSYS_UNCONNECTED_945, 
        SYNOPSYS_UNCONNECTED_946, SYNOPSYS_UNCONNECTED_947, 
        SYNOPSYS_UNCONNECTED_948, SYNOPSYS_UNCONNECTED_949, 
        SYNOPSYS_UNCONNECTED_950, SYNOPSYS_UNCONNECTED_951, 
        SYNOPSYS_UNCONNECTED_952, SYNOPSYS_UNCONNECTED_953, 
        SYNOPSYS_UNCONNECTED_954, SYNOPSYS_UNCONNECTED_955, 
        SYNOPSYS_UNCONNECTED_956, SYNOPSYS_UNCONNECTED_957, 
        SYNOPSYS_UNCONNECTED_958, SYNOPSYS_UNCONNECTED_959, 
        SYNOPSYS_UNCONNECTED_960, SYNOPSYS_UNCONNECTED_961, 
        SYNOPSYS_UNCONNECTED_962, SYNOPSYS_UNCONNECTED_963, 
        SYNOPSYS_UNCONNECTED_964, SYNOPSYS_UNCONNECTED_965, 
        SYNOPSYS_UNCONNECTED_966, SYNOPSYS_UNCONNECTED_967, 
        SYNOPSYS_UNCONNECTED_968, SYNOPSYS_UNCONNECTED_969, 
        SYNOPSYS_UNCONNECTED_970, SYNOPSYS_UNCONNECTED_971, 
        SYNOPSYS_UNCONNECTED_972, SYNOPSYS_UNCONNECTED_973, 
        SYNOPSYS_UNCONNECTED_974, SYNOPSYS_UNCONNECTED_975, 
        SYNOPSYS_UNCONNECTED_976, SYNOPSYS_UNCONNECTED_977, 
        SYNOPSYS_UNCONNECTED_978, SYNOPSYS_UNCONNECTED_979, 
        SYNOPSYS_UNCONNECTED_980, SYNOPSYS_UNCONNECTED_981, 
        SYNOPSYS_UNCONNECTED_982, SYNOPSYS_UNCONNECTED_983, 
        SYNOPSYS_UNCONNECTED_984, SYNOPSYS_UNCONNECTED_985, 
        SYNOPSYS_UNCONNECTED_986, SYNOPSYS_UNCONNECTED_987, 
        SYNOPSYS_UNCONNECTED_988, SYNOPSYS_UNCONNECTED_989, 
        SYNOPSYS_UNCONNECTED_990, SYNOPSYS_UNCONNECTED_991, 
        SYNOPSYS_UNCONNECTED_992, SYNOPSYS_UNCONNECTED_993, 
        SYNOPSYS_UNCONNECTED_994, SYNOPSYS_UNCONNECTED_995, 
        SYNOPSYS_UNCONNECTED_996, SYNOPSYS_UNCONNECTED_997, 
        SYNOPSYS_UNCONNECTED_998, SYNOPSYS_UNCONNECTED_999, 
        SYNOPSYS_UNCONNECTED_1000, SYNOPSYS_UNCONNECTED_1001, 
        SYNOPSYS_UNCONNECTED_1002, SYNOPSYS_UNCONNECTED_1003, 
        SYNOPSYS_UNCONNECTED_1004, SYNOPSYS_UNCONNECTED_1005, 
        SYNOPSYS_UNCONNECTED_1006, SYNOPSYS_UNCONNECTED_1007, 
        SYNOPSYS_UNCONNECTED_1008, SYNOPSYS_UNCONNECTED_1009, 
        SYNOPSYS_UNCONNECTED_1010, SYNOPSYS_UNCONNECTED_1011, 
        SYNOPSYS_UNCONNECTED_1012, SYNOPSYS_UNCONNECTED_1013, 
        SYNOPSYS_UNCONNECTED_1014, SYNOPSYS_UNCONNECTED_1015, 
        SYNOPSYS_UNCONNECTED_1016, SYNOPSYS_UNCONNECTED_1017, sfr_rdat}) );
  HAD1X1 add_179_U1_1_1 ( .A(N26), .B(N27), .CO(add_179_carry[2]), .SO(N29) );
  HAD1X1 add_179_U1_1_2 ( .A(N25), .B(add_179_carry[2]), .CO(add_179_carry[3]), 
        .SO(N30) );
  HAD1X1 add_179_U1_1_3 ( .A(N24), .B(add_179_carry[3]), .CO(add_179_carry[4]), 
        .SO(N31) );
  DFFRQX1 r_phyrst_reg_0_ ( .D(n1210), .C(clk), .XR(n6), .Q(r_phyrst[0]) );
  DFFRQX1 rstcnt_reg_0_ ( .D(N36), .C(net10758), .XR(n7), .Q(rstcnt[0]) );
  DFFRQX1 d_p0_reg_7_ ( .D(ff_p0[7]), .C(clk), .XR(n294), .Q(d_p0[7]) );
  DFFRQX1 d_p0_reg_6_ ( .D(ff_p0[6]), .C(clk), .XR(n294), .Q(d_p0[6]) );
  DFFRQX1 d_p0_reg_5_ ( .D(ff_p0[5]), .C(clk), .XR(n294), .Q(d_p0[5]) );
  DFFRQX1 d_p0_reg_4_ ( .D(ff_p0[4]), .C(clk), .XR(n294), .Q(d_p0[4]) );
  DFFRQX1 d_p0_reg_3_ ( .D(ff_p0[3]), .C(clk), .XR(n294), .Q(d_p0[3]) );
  DFFRQX1 d_p0_reg_2_ ( .D(ff_p0[2]), .C(clk), .XR(n294), .Q(d_p0[2]) );
  DFFRQX1 d_p0_reg_1_ ( .D(ff_p0[1]), .C(clk), .XR(n294), .Q(d_p0[1]) );
  DFFRQX1 d_p0_reg_0_ ( .D(ff_p0[0]), .C(clk), .XR(n294), .Q(d_p0[0]) );
  DFFRQX1 r_phyrst_reg_1_ ( .D(n1209), .C(clk), .XR(n6), .Q(r_phyrst[1]) );
  DFFQX1 oscdwn_shft_reg_2_ ( .D(n238), .C(clk), .Q(oscdwn_shft[2]) );
  DFFQX1 oscdwn_shft_reg_1_ ( .D(oscdwn_shft[0]), .C(clk), .Q(oscdwn_shft[1])
         );
  DFFNRQX1 osc_gate_n_reg_3_ ( .D(osc_gate_n[2]), .XC(xclk), .XR(n6), .Q(
        osc_gate_n[3]) );
  DFFNRQX1 osc_gate_n_reg_0_ ( .D(r_pos_gate), .XC(xclk), .XR(n7), .Q(
        osc_gate_n[0]) );
  DFFNRQX1 osc_gate_n_reg_1_ ( .D(osc_gate_n[0]), .XC(xclk), .XR(n7), .Q(
        osc_gate_n[1]) );
  DFFNRQX1 osc_gate_n_reg_2_ ( .D(osc_gate_n[1]), .XC(xclk), .XR(n6), .Q(
        osc_gate_n[2]) );
  DFFRQX1 rstcnt_reg_1_ ( .D(N35), .C(net10758), .XR(n7), .Q(rstcnt[1]) );
  DFFRQX1 rstcnt_reg_2_ ( .D(N34), .C(net10758), .XR(n6), .Q(rstcnt[2]) );
  DFFRQX1 drstz_reg_1_ ( .D(drstz[0]), .C(clk), .XR(n6), .Q(drstz[1]) );
  DFFRQX1 rstcnt_reg_4_ ( .D(N32), .C(net10758), .XR(n7), .Q(rstcnt[4]) );
  DFFRQX1 rstcnt_reg_3_ ( .D(N33), .C(net10758), .XR(n6), .Q(rstcnt[3]) );
  DFFQX1 oscdwn_shft_reg_0_ ( .D(N81), .C(clk), .Q(oscdwn_shft[0]) );
  DFFRQX1 drstz_reg_0_ ( .D(1'b1), .C(clk), .XR(n7), .Q(drstz[0]) );
  NAND21X1 U3 ( .B(n206), .A(sfr_addr[2]), .Y(n226) );
  NOR2X1 U4 ( .A(n216), .B(n240), .Y(n31) );
  INVX1 U5 ( .A(n225), .Y(n4) );
  INVX1 U6 ( .A(n225), .Y(n274) );
  NAND21X1 U10 ( .B(n258), .A(n224), .Y(n225) );
  INVX1 U11 ( .A(xrstz), .Y(n5) );
  INVX1 U12 ( .A(n5), .Y(n6) );
  INVX1 U13 ( .A(n5), .Y(n7) );
  INVX1 U14 ( .A(n253), .Y(n8) );
  INVX1 U15 ( .A(n227), .Y(n9) );
  BUFX3 U16 ( .A(n1125), .Y(n10) );
  INVX1 U17 ( .A(n1133), .Y(n11) );
  INVX1 U18 ( .A(n219), .Y(n12) );
  INVX1 U19 ( .A(n280), .Y(n13) );
  BUFX3 U20 ( .A(n275), .Y(n14) );
  AND2X1 U21 ( .A(pff_ack[0]), .B(n14), .Y(set04[4]) );
  BUFX3 U22 ( .A(n1126), .Y(n15) );
  NAND21X1 U23 ( .B(n223), .A(n71), .Y(n258) );
  BUFX3 U24 ( .A(phyrst), .Y(n16) );
  BUFX3 U25 ( .A(pff_ptr[4]), .Y(dbgpo[20]) );
  BUFX3 U26 ( .A(pff_ptr[0]), .Y(dbgpo[16]) );
  BUFX3 U27 ( .A(pff_ptr[2]), .Y(dbgpo[18]) );
  BUFX3 U28 ( .A(pff_ptr[1]), .Y(dbgpo[17]) );
  BUFX3 U29 ( .A(pff_ptr[3]), .Y(dbgpo[19]) );
  BUFX3 U30 ( .A(pff_ptr[5]), .Y(dbgpo[21]) );
  NAND21XL U31 ( .B(n221), .A(n220), .Y(n222) );
  NAND32XL U32 ( .B(n245), .C(n221), .A(n152), .Y(n207) );
  NAND32XL U33 ( .B(n245), .C(n152), .A(n244), .Y(n228) );
  NAND32XL U34 ( .B(n245), .C(n244), .A(n152), .Y(n246) );
  NAND21XL U35 ( .B(n244), .A(n220), .Y(n253) );
  NAND21X1 U36 ( .B(n206), .A(sfr_addr[4]), .Y(n240) );
  NAND21XL U37 ( .B(n76), .A(n224), .Y(n218) );
  NOR2XL U38 ( .A(n242), .B(n216), .Y(n62) );
  NAND21XL U39 ( .B(n242), .A(n241), .Y(n204) );
  NAND21XL U40 ( .B(n242), .A(n239), .Y(n212) );
  INVXL U41 ( .A(sfr_addr[6]), .Y(n156) );
  NAND31X1 U42 ( .C(n240), .A(n302), .B(n236), .Y(n213) );
  NAND21XL U43 ( .B(n206), .A(sfr_addr[1]), .Y(n244) );
  NAND21XL U44 ( .B(n206), .A(sfr_addr[3]), .Y(n236) );
  ENOXL U45 ( .A(n161), .B(n1136), .C(r_txnumk[0]), .D(n1136), .Y(wd01[0]) );
  ENOXL U46 ( .A(n167), .B(n13), .C(r_txnumk[1]), .D(n1136), .Y(wd01[1]) );
  ENOXL U47 ( .A(n173), .B(n13), .C(r_txnumk[2]), .D(n1136), .Y(wd01[2]) );
  ENOXL U48 ( .A(n178), .B(n13), .C(r_txnumk[3]), .D(n1136), .Y(wd01[3]) );
  INVX3 U49 ( .A(n157), .Y(n155) );
  INVX1 U50 ( .A(n179), .Y(n174) );
  INVX1 U51 ( .A(n72), .Y(n74) );
  INVX1 U52 ( .A(n71), .Y(n75) );
  INVX1 U53 ( .A(n72), .Y(n76) );
  NAND4XL U54 ( .A(n279), .B(n174), .C(n1177), .D(n191), .Y(n1149) );
  NOR2X1 U55 ( .A(n160), .B(n201), .Y(n1177) );
  NOR3XL U56 ( .A(n1149), .B(n185), .C(n173), .Y(r_discard) );
  INVX1 U57 ( .A(n218), .Y(n229) );
  INVX1 U58 ( .A(n195), .Y(n191) );
  INVX1 U59 ( .A(n72), .Y(n73) );
  INVX1 U60 ( .A(n172), .Y(n168) );
  INVX1 U61 ( .A(n202), .Y(n197) );
  INVX1 U62 ( .A(n195), .Y(n194) );
  INVX1 U63 ( .A(n201), .Y(n200) );
  INVX1 U64 ( .A(n184), .Y(n182) );
  INVX1 U65 ( .A(n201), .Y(n199) );
  INVX1 U66 ( .A(n161), .Y(n159) );
  INVX1 U67 ( .A(n167), .Y(n164) );
  INVX1 U68 ( .A(n190), .Y(n187) );
  INVX1 U69 ( .A(n196), .Y(n193) );
  INVX1 U70 ( .A(n173), .Y(n170) );
  INVX1 U71 ( .A(n178), .Y(n175) );
  INVX1 U72 ( .A(n195), .Y(n192) );
  INVX1 U73 ( .A(n201), .Y(n198) );
  INVX1 U74 ( .A(n161), .Y(n158) );
  INVX1 U75 ( .A(n173), .Y(n169) );
  INVX1 U76 ( .A(n190), .Y(n186) );
  INVX1 U77 ( .A(n166), .Y(n163) );
  INVX1 U78 ( .A(n184), .Y(n181) );
  INVX1 U79 ( .A(n178), .Y(n176) );
  INVX1 U80 ( .A(n184), .Y(n180) );
  INVX1 U81 ( .A(n190), .Y(n188) );
  INVX1 U82 ( .A(n185), .Y(n183) );
  INVX1 U83 ( .A(n172), .Y(n171) );
  INVX1 U84 ( .A(n162), .Y(n160) );
  INVX1 U85 ( .A(n166), .Y(n165) );
  INVX1 U86 ( .A(n178), .Y(n177) );
  INVX1 U87 ( .A(n135), .Y(n129) );
  INVX1 U88 ( .A(n139), .Y(n128) );
  INVX1 U89 ( .A(n145), .Y(n127) );
  INVX1 U90 ( .A(n147), .Y(n84) );
  INVX1 U91 ( .A(n135), .Y(n130) );
  INVX1 U92 ( .A(n148), .Y(n133) );
  INVX1 U93 ( .A(n142), .Y(n132) );
  INVX1 U94 ( .A(n140), .Y(n96) );
  INVX1 U95 ( .A(n138), .Y(n117) );
  INVX1 U96 ( .A(n138), .Y(n119) );
  INVX1 U97 ( .A(n148), .Y(n86) );
  INVX1 U98 ( .A(n143), .Y(n92) );
  INVX1 U99 ( .A(n147), .Y(n94) );
  INVX1 U100 ( .A(n136), .Y(n89) );
  INVX1 U101 ( .A(n143), .Y(n90) );
  INVX1 U102 ( .A(n143), .Y(n91) );
  INVX1 U103 ( .A(n139), .Y(n98) );
  INVX1 U104 ( .A(n147), .Y(n102) );
  INVX1 U105 ( .A(n144), .Y(n95) );
  INVX1 U106 ( .A(n135), .Y(n131) );
  INVX1 U107 ( .A(n145), .Y(n104) );
  INVX1 U108 ( .A(n141), .Y(n105) );
  INVX1 U109 ( .A(n140), .Y(n110) );
  INVX1 U110 ( .A(n141), .Y(n107) );
  INVX1 U111 ( .A(n140), .Y(n108) );
  INVX1 U112 ( .A(n140), .Y(n109) );
  INVX1 U113 ( .A(n139), .Y(n114) );
  INVX1 U114 ( .A(n142), .Y(n111) );
  INVX1 U115 ( .A(n147), .Y(n113) );
  INVX1 U116 ( .A(n139), .Y(n115) );
  INVX1 U117 ( .A(n139), .Y(n116) );
  INVX1 U118 ( .A(n138), .Y(n118) );
  INVX1 U119 ( .A(n137), .Y(n120) );
  INVX1 U120 ( .A(n1211), .Y(n112) );
  INVX1 U121 ( .A(n141), .Y(n106) );
  INVX1 U122 ( .A(n142), .Y(n101) );
  INVX1 U123 ( .A(n142), .Y(n100) );
  INVX1 U124 ( .A(n142), .Y(n99) );
  INVX1 U125 ( .A(n138), .Y(n97) );
  INVX1 U126 ( .A(n143), .Y(n93) );
  INVX1 U127 ( .A(n137), .Y(n88) );
  INVX1 U128 ( .A(n148), .Y(n87) );
  INVX1 U129 ( .A(n141), .Y(n85) );
  INVX1 U130 ( .A(n135), .Y(n103) );
  INVX1 U131 ( .A(n137), .Y(n121) );
  INVX1 U132 ( .A(n137), .Y(n122) );
  INVX1 U133 ( .A(n136), .Y(n123) );
  INVX1 U134 ( .A(n136), .Y(n124) );
  INVX1 U135 ( .A(n136), .Y(n125) );
  INVX1 U136 ( .A(n135), .Y(n126) );
  INVX1 U137 ( .A(n144), .Y(n134) );
  INVX1 U138 ( .A(atpg_en), .Y(n203) );
  INVX1 U139 ( .A(n217), .Y(n224) );
  INVX1 U140 ( .A(sfr_wdat[3]), .Y(n179) );
  NOR2X1 U141 ( .A(n17), .B(n75), .Y(r_dacwr[7]) );
  NAND2X1 U142 ( .A(n248), .B(n8), .Y(n17) );
  NOR2X1 U143 ( .A(n18), .B(n75), .Y(r_dacwr[5]) );
  NAND2X1 U144 ( .A(n248), .B(n271), .Y(n18) );
  AND2X1 U145 ( .A(n34), .B(n248), .Y(r_dacwr[4]) );
  NOR2X1 U146 ( .A(n19), .B(n76), .Y(r_dacwr[0]) );
  NAND2X1 U147 ( .A(n248), .B(n263), .Y(n19) );
  INVX1 U148 ( .A(sfr_wdat[7]), .Y(n201) );
  INVX1 U149 ( .A(sfr_wdat[6]), .Y(n195) );
  INVX1 U150 ( .A(sfr_wdat[0]), .Y(n161) );
  INVX1 U151 ( .A(sfr_wdat[2]), .Y(n172) );
  INVX1 U152 ( .A(sfr_wdat[4]), .Y(n184) );
  INVX1 U153 ( .A(sfr_wdat[3]), .Y(n178) );
  INVX1 U154 ( .A(sfr_wdat[1]), .Y(n166) );
  INVX1 U155 ( .A(sfr_wdat[5]), .Y(n189) );
  AND2X1 U156 ( .A(n34), .B(n249), .Y(r_fcpwr[1]) );
  NOR2X1 U157 ( .A(n202), .B(n1124), .Y(r_i2c_fwack) );
  NOR2X1 U158 ( .A(n20), .B(n74), .Y(r_fcpwr[5]) );
  NAND2X1 U159 ( .A(n249), .B(n269), .Y(n20) );
  AND2X1 U160 ( .A(n34), .B(n272), .Y(r_dacwr[11]) );
  NOR2X1 U161 ( .A(n189), .B(n1185), .Y(clr28[5]) );
  NOR2X1 U162 ( .A(n167), .B(n1185), .Y(clr28[1]) );
  NOR2X1 U163 ( .A(n189), .B(n1186), .Y(clr04[5]) );
  NOR2X1 U164 ( .A(n167), .B(n1186), .Y(clr04[1]) );
  NOR2X1 U165 ( .A(n185), .B(n1185), .Y(clr28[4]) );
  NOR2X1 U166 ( .A(n162), .B(n1185), .Y(clr28[0]) );
  NOR2X1 U167 ( .A(n185), .B(n1186), .Y(clr04[4]) );
  NOR2X1 U168 ( .A(n162), .B(n1186), .Y(clr04[0]) );
  NOR2X1 U169 ( .A(n196), .B(n1124), .Y(r_i2c_fwnak) );
  INVX1 U170 ( .A(n1147), .Y(n279) );
  NOR2X1 U171 ( .A(n21), .B(n74), .Y(r_pwrv_upd) );
  NAND2X1 U172 ( .A(n270), .B(n271), .Y(n21) );
  AND3X1 U173 ( .A(n215), .B(n302), .C(n269), .Y(we_143) );
  AND2X1 U174 ( .A(n34), .B(n270), .Y(we_228) );
  AND2X1 U175 ( .A(n34), .B(n262), .Y(we_172) );
  AND2X1 U176 ( .A(n229), .B(n269), .Y(we_215) );
  AND2X1 U177 ( .A(n229), .B(n271), .Y(we_213) );
  AND2X1 U178 ( .A(n34), .B(n261), .Y(we[164]) );
  NOR2X1 U179 ( .A(n196), .B(n1185), .Y(clr28[6]) );
  NOR2X1 U180 ( .A(n173), .B(n1185), .Y(clr28[2]) );
  NOR2X1 U181 ( .A(n196), .B(n1186), .Y(clr04[6]) );
  NOR2X1 U182 ( .A(n172), .B(n1186), .Y(clr04[2]) );
  NOR2X1 U183 ( .A(n202), .B(n1185), .Y(clr28[7]) );
  NOR2X1 U184 ( .A(n178), .B(n1185), .Y(clr28[3]) );
  NOR2X1 U185 ( .A(n202), .B(n1186), .Y(clr04[7]) );
  NOR2X1 U186 ( .A(n178), .B(n1186), .Y(clr04[3]) );
  INVX1 U187 ( .A(sfr_wdat[0]), .Y(n162) );
  NOR2X1 U188 ( .A(n189), .B(n1184), .Y(clrAE[5]) );
  NOR2X1 U189 ( .A(n167), .B(n1184), .Y(clrAE[1]) );
  NOR2X1 U190 ( .A(n189), .B(n1183), .Y(clrDF[5]) );
  NOR2X1 U191 ( .A(n166), .B(n1183), .Y(clrDF[1]) );
  NOR2X1 U192 ( .A(n189), .B(n1187), .Y(clr03[5]) );
  NOR2X1 U193 ( .A(n167), .B(n1187), .Y(clr03[1]) );
  NOR2X1 U194 ( .A(n184), .B(n1184), .Y(clrAE[4]) );
  NOR2X1 U195 ( .A(n162), .B(n1184), .Y(clrAE[0]) );
  NOR2X1 U196 ( .A(n185), .B(n1183), .Y(clrDF[4]) );
  NOR2X1 U197 ( .A(n162), .B(n1183), .Y(clrDF[0]) );
  NOR2X1 U198 ( .A(n184), .B(n1187), .Y(clr03[4]) );
  NOR2X1 U199 ( .A(n162), .B(n1187), .Y(clr03[0]) );
  NOR2X1 U200 ( .A(n196), .B(n1184), .Y(clrAE[6]) );
  NOR2X1 U201 ( .A(n173), .B(n1184), .Y(clrAE[2]) );
  NOR2X1 U202 ( .A(n196), .B(n1183), .Y(clrDF[6]) );
  NOR2X1 U203 ( .A(n172), .B(n1183), .Y(clrDF[2]) );
  NOR2X1 U204 ( .A(n196), .B(n1187), .Y(clr03[6]) );
  NOR2X1 U205 ( .A(n173), .B(n1187), .Y(clr03[2]) );
  NOR2X1 U206 ( .A(n202), .B(n1184), .Y(clrAE[7]) );
  NOR2X1 U207 ( .A(n178), .B(n1184), .Y(clrAE[3]) );
  NOR2X1 U208 ( .A(n202), .B(n1183), .Y(clrDF[7]) );
  NOR2X1 U209 ( .A(n178), .B(n1183), .Y(clrDF[3]) );
  NOR2X1 U210 ( .A(n202), .B(n1187), .Y(clr03[7]) );
  NOR2X1 U211 ( .A(n178), .B(n1187), .Y(clr03[3]) );
  INVX1 U212 ( .A(n205), .Y(n215) );
  NAND21X1 U213 ( .B(n76), .A(n209), .Y(n205) );
  INVX1 U214 ( .A(n257), .Y(n259) );
  NAND21X1 U215 ( .B(n1128), .A(n151), .Y(n1127) );
  NOR2X1 U216 ( .A(n22), .B(n74), .Y(r_fcpwr[2]) );
  NAND2X1 U217 ( .A(n249), .B(n271), .Y(n22) );
  NOR2X1 U218 ( .A(n23), .B(n73), .Y(we_245) );
  NAND2X1 U219 ( .A(n271), .B(n272), .Y(n23) );
  NOR2X1 U220 ( .A(n24), .B(n73), .Y(we_231) );
  NAND2X1 U221 ( .A(n270), .B(n269), .Y(n24) );
  NOR2X1 U222 ( .A(n25), .B(n76), .Y(we_175) );
  NAND2X1 U223 ( .A(n262), .B(n269), .Y(n25) );
  NOR2X1 U224 ( .A(n26), .B(n76), .Y(we[167]) );
  NAND2X1 U225 ( .A(n261), .B(n269), .Y(n26) );
  NOR2X1 U226 ( .A(n27), .B(n76), .Y(we[165]) );
  NAND2X1 U227 ( .A(n261), .B(n271), .Y(n27) );
  NOR2X1 U228 ( .A(n28), .B(n73), .Y(we_191) );
  NAND2X1 U229 ( .A(n265), .B(n269), .Y(n28) );
  NOR2X1 U230 ( .A(n29), .B(n76), .Y(we_181) );
  NAND2X1 U231 ( .A(n264), .B(n271), .Y(n29) );
  NOR2X1 U232 ( .A(n30), .B(n277), .Y(we_176) );
  NAND2X1 U233 ( .A(n263), .B(n264), .Y(n30) );
  INVX1 U234 ( .A(sfr_wdat[2]), .Y(n173) );
  INVX1 U235 ( .A(sfr_wdat[4]), .Y(n185) );
  INVX1 U236 ( .A(sfr_wdat[6]), .Y(n196) );
  INVX1 U237 ( .A(sfr_wdat[7]), .Y(n202) );
  INVX1 U238 ( .A(n1136), .Y(n280) );
  INVX1 U239 ( .A(n1123), .Y(n1095) );
  INVX1 U240 ( .A(n1124), .Y(n1096) );
  INVX1 U241 ( .A(sfr_wdat[5]), .Y(n190) );
  INVX1 U242 ( .A(sfr_wdat[1]), .Y(n167) );
  INVX1 U243 ( .A(n151), .Y(n149) );
  INVX1 U244 ( .A(n151), .Y(n150) );
  INVX1 U245 ( .A(n145), .Y(n78) );
  INVX1 U246 ( .A(n145), .Y(n79) );
  INVX1 U247 ( .A(n145), .Y(n80) );
  INVX1 U248 ( .A(n144), .Y(n81) );
  INVX1 U249 ( .A(n144), .Y(n82) );
  INVX1 U250 ( .A(n144), .Y(n83) );
  INVX1 U251 ( .A(n146), .Y(n143) );
  INVX1 U252 ( .A(n146), .Y(n136) );
  INVX1 U253 ( .A(n1076), .Y(n135) );
  INVX1 U254 ( .A(n1076), .Y(n139) );
  INVX1 U255 ( .A(n146), .Y(n138) );
  INVX1 U256 ( .A(n146), .Y(n137) );
  INVX1 U257 ( .A(n146), .Y(n141) );
  INVX1 U258 ( .A(n1076), .Y(n142) );
  INVX1 U259 ( .A(n146), .Y(n140) );
  NAND21X1 U260 ( .B(n241), .A(n155), .Y(n216) );
  INVX1 U261 ( .A(n154), .Y(n153) );
  INVX1 U262 ( .A(sfr_addr[0]), .Y(n152) );
  NOR2X1 U263 ( .A(n32), .B(n74), .Y(r_dacwr[8]) );
  NAND2X1 U264 ( .A(n267), .B(n272), .Y(n32) );
  INVX1 U265 ( .A(n72), .Y(n277) );
  NOR2X1 U266 ( .A(n33), .B(n75), .Y(r_dacwr[6]) );
  NAND2X1 U267 ( .A(n248), .B(n273), .Y(n33) );
  NOR2X1 U268 ( .A(n76), .B(n223), .Y(n34) );
  NOR2X1 U269 ( .A(n35), .B(n75), .Y(r_dacwr[2]) );
  NAND2X1 U270 ( .A(n248), .B(n260), .Y(n35) );
  NOR2X1 U271 ( .A(n36), .B(n75), .Y(r_dacwr[1]) );
  NAND2X1 U272 ( .A(n248), .B(n267), .Y(n36) );
  NOR2X1 U273 ( .A(n37), .B(n75), .Y(r_dacwr[3]) );
  NAND2X1 U274 ( .A(n248), .B(n9), .Y(n37) );
  OAI31XL U275 ( .A(n1146), .B(n1147), .C(n1148), .D(n284), .Y(r_fiforst) );
  NAND2X1 U276 ( .A(n161), .B(n172), .Y(n1148) );
  NAND4X1 U277 ( .A(n178), .B(n184), .C(n195), .D(n201), .Y(n1146) );
  INVX1 U278 ( .A(n233), .Y(n248) );
  INVX1 U279 ( .A(n234), .Y(n272) );
  NAND4X1 U280 ( .A(hit[183]), .B(n71), .C(n166), .D(n189), .Y(n1147) );
  AND2X1 U281 ( .A(n264), .B(n269), .Y(hit[183]) );
  INVX1 U282 ( .A(n253), .Y(n269) );
  INVX1 U283 ( .A(n222), .Y(n271) );
  INVX1 U284 ( .A(n207), .Y(n263) );
  NOR2X1 U285 ( .A(n38), .B(n74), .Y(r_fcpwr[3]) );
  NAND2X1 U286 ( .A(n249), .B(n273), .Y(n38) );
  INVX1 U287 ( .A(n211), .Y(n239) );
  INVX1 U288 ( .A(n243), .Y(n266) );
  INVX1 U289 ( .A(n251), .Y(n264) );
  AND2X1 U290 ( .A(hit[178]), .B(n72), .Y(r_fifopsh) );
  INVX1 U291 ( .A(n254), .Y(hit_207) );
  NAND21X1 U292 ( .B(n253), .A(n266), .Y(n254) );
  INVX1 U293 ( .A(n252), .Y(hit[178]) );
  NAND21X1 U294 ( .B(n251), .A(n260), .Y(n252) );
  NOR2X1 U295 ( .A(n39), .B(n75), .Y(r_dacwr[12]) );
  NAND2X1 U296 ( .A(n260), .B(n270), .Y(n39) );
  INVX1 U297 ( .A(n235), .Y(n249) );
  NAND21X1 U298 ( .B(n255), .A(n302), .Y(n235) );
  NOR2X1 U299 ( .A(n40), .B(n74), .Y(r_fcpwr[4]) );
  NAND2X1 U300 ( .A(n250), .B(n271), .Y(n40) );
  NAND2X1 U301 ( .A(hit_201), .B(n72), .Y(n1124) );
  AND2X1 U302 ( .A(n266), .B(n267), .Y(hit_201) );
  NOR2X1 U303 ( .A(n41), .B(n74), .Y(r_set_cpmsgid) );
  NAND2X1 U304 ( .A(n265), .B(n273), .Y(n41) );
  NAND2X1 U305 ( .A(hit[174]), .B(n71), .Y(n1184) );
  AND2X1 U306 ( .A(n262), .B(n273), .Y(hit[174]) );
  NAND2X1 U307 ( .A(hit_223), .B(n72), .Y(n1183) );
  AND2X1 U308 ( .A(n43), .B(n269), .Y(hit_223) );
  NAND2X1 U309 ( .A(hit[179]), .B(n71), .Y(n1187) );
  AND2X1 U310 ( .A(n264), .B(n268), .Y(hit[179]) );
  NAND2X1 U311 ( .A(hit_202), .B(n72), .Y(n1123) );
  AND2X1 U312 ( .A(n260), .B(n266), .Y(hit_202) );
  AND2X1 U313 ( .A(n229), .B(n12), .Y(we_214) );
  AND2X1 U314 ( .A(n34), .B(n247), .Y(r_cvcwr[0]) );
  AND2X1 U315 ( .A(n229), .B(n268), .Y(we_211) );
  AND2X1 U316 ( .A(n229), .B(n267), .Y(we_209) );
  AND2X1 U317 ( .A(n34), .B(n250), .Y(we_148) );
  INVX1 U318 ( .A(prl_c0set), .Y(n284) );
  NAND2X1 U319 ( .A(hit[177]), .B(n71), .Y(n1136) );
  AND2X1 U320 ( .A(n264), .B(n267), .Y(hit[177]) );
  AND2X1 U321 ( .A(n259), .B(n260), .Y(hit_194) );
  INVX1 U322 ( .A(n204), .Y(n209) );
  NAND2X1 U323 ( .A(hit_197), .B(n72), .Y(n1125) );
  AND2X1 U324 ( .A(n259), .B(n271), .Y(hit_197) );
  NOR2X1 U325 ( .A(n42), .B(n76), .Y(we[162]) );
  NAND2X1 U326 ( .A(n260), .B(n261), .Y(n42) );
  NOR3XL U327 ( .A(n156), .B(n153), .C(n255), .Y(n43) );
  INVX1 U328 ( .A(n210), .Y(n262) );
  NOR2X1 U329 ( .A(n44), .B(n74), .Y(r_fcpwr[0]) );
  NAND2X1 U330 ( .A(n249), .B(n268), .Y(n44) );
  NOR2X1 U331 ( .A(n45), .B(n74), .Y(r_fcpwr[6]) );
  NAND2X1 U332 ( .A(n250), .B(n273), .Y(n45) );
  NOR2X1 U333 ( .A(n46), .B(n76), .Y(r_cvcwr[1]) );
  NAND2X1 U334 ( .A(n247), .B(n271), .Y(n46) );
  NOR2X1 U335 ( .A(n47), .B(n75), .Y(r_dacwr[14]) );
  NAND2X1 U336 ( .A(n250), .B(n267), .Y(n47) );
  NOR2X1 U337 ( .A(n48), .B(n75), .Y(r_dacwr[13]) );
  NAND2X1 U338 ( .A(n250), .B(n263), .Y(n48) );
  NOR2X1 U339 ( .A(n49), .B(n75), .Y(r_dacwr[10]) );
  NAND2X1 U340 ( .A(n268), .B(n272), .Y(n49) );
  NOR2X1 U341 ( .A(n50), .B(n74), .Y(r_dacwr[9]) );
  NAND2X1 U342 ( .A(n260), .B(n272), .Y(n50) );
  NOR2X1 U343 ( .A(n51), .B(n73), .Y(we_246) );
  NAND2X1 U344 ( .A(n12), .B(n272), .Y(n51) );
  NOR2X1 U345 ( .A(n52), .B(n73), .Y(we_230) );
  NAND2X1 U346 ( .A(n270), .B(n273), .Y(n52) );
  NOR2X1 U347 ( .A(n53), .B(n73), .Y(we_227) );
  NAND2X1 U348 ( .A(n268), .B(n270), .Y(n53) );
  NOR2X1 U349 ( .A(n54), .B(n277), .Y(we_171) );
  NAND2X1 U350 ( .A(n262), .B(n268), .Y(n54) );
  NOR2X1 U351 ( .A(n55), .B(n277), .Y(we[166]) );
  NAND2X1 U352 ( .A(n261), .B(n273), .Y(n55) );
  NOR2X1 U353 ( .A(n56), .B(n277), .Y(we[163]) );
  NAND2X1 U354 ( .A(n261), .B(n268), .Y(n56) );
  NOR2X1 U355 ( .A(n57), .B(n73), .Y(we_222) );
  NAND2X1 U356 ( .A(n43), .B(n273), .Y(n57) );
  NOR2X1 U357 ( .A(n58), .B(n73), .Y(we_217) );
  NAND2X1 U358 ( .A(n267), .B(n43), .Y(n58) );
  NOR2X1 U359 ( .A(n59), .B(n73), .Y(we_203) );
  NAND2X1 U360 ( .A(n266), .B(n268), .Y(n59) );
  NOR2X1 U361 ( .A(n60), .B(n73), .Y(we_187) );
  NAND2X1 U362 ( .A(n265), .B(n268), .Y(n60) );
  NOR2X1 U363 ( .A(n61), .B(n277), .Y(we_182) );
  NAND2X1 U364 ( .A(n264), .B(n273), .Y(n61) );
  NAND2X1 U365 ( .A(hit_195), .B(n71), .Y(n1128) );
  AND2X1 U366 ( .A(n259), .B(n268), .Y(hit_195) );
  INVX1 U367 ( .A(n1133), .Y(n281) );
  INVX1 U368 ( .A(n208), .Y(n270) );
  INVX1 U369 ( .A(n256), .Y(n265) );
  INVX1 U370 ( .A(n212), .Y(n261) );
  INVX1 U371 ( .A(ictlr_inc), .Y(n151) );
  INVX1 U372 ( .A(n148), .Y(n77) );
  INVX1 U373 ( .A(n148), .Y(n146) );
  INVX1 U374 ( .A(n1076), .Y(n145) );
  INVX1 U375 ( .A(n1076), .Y(n144) );
  NAND32X1 U376 ( .B(n221), .C(n226), .A(n152), .Y(n223) );
  INVX1 U377 ( .A(n236), .Y(n241) );
  INVX1 U378 ( .A(n240), .Y(n242) );
  INVX1 U379 ( .A(n244), .Y(n221) );
  INVX1 U380 ( .A(sfr_addr[6]), .Y(n157) );
  NAND21XL U381 ( .B(n240), .A(n241), .Y(n255) );
  INVX1 U382 ( .A(n228), .Y(n267) );
  INVX1 U383 ( .A(n214), .Y(n220) );
  NAND21XL U384 ( .B(n226), .A(sfr_addr[0]), .Y(n214) );
  INVXL U385 ( .A(n226), .Y(n245) );
  INVX1 U386 ( .A(n219), .Y(n273) );
  NAND32XL U387 ( .B(n244), .C(n226), .A(n152), .Y(n219) );
  INVX1 U388 ( .A(n227), .Y(n268) );
  NAND32XL U389 ( .B(n244), .C(n152), .A(n226), .Y(n227) );
  NAND21X1 U390 ( .B(n240), .A(n239), .Y(n251) );
  AND2X1 U391 ( .A(sfr_r), .B(hit[178]), .Y(r_fifopop) );
  INVX1 U392 ( .A(n246), .Y(n260) );
  OA21X1 U393 ( .B(prx_rst[0]), .C(prx_rst[1]), .A(set03[1]), .Y(set03[7]) );
  AND2X1 U394 ( .A(hit_151), .B(sfr_r), .Y(r_fcpre) );
  AND2X1 U395 ( .A(n250), .B(n269), .Y(hit_151) );
  INVX1 U396 ( .A(n1152), .Y(n278) );
  NOR2X1 U397 ( .A(n1129), .B(n296), .Y(n1133) );
  NAND4X1 U398 ( .A(n1128), .B(n278), .C(n1141), .D(n151), .Y(upd19) );
  INVX1 U399 ( .A(n213), .Y(n250) );
  INVX1 U400 ( .A(n237), .Y(n247) );
  INVX1 U401 ( .A(n1140), .Y(n1120) );
  INVX1 U402 ( .A(N31), .Y(n297) );
  INVX1 U403 ( .A(n1076), .Y(n147) );
  INVX1 U404 ( .A(n1076), .Y(n148) );
  BUFX3 U405 ( .A(pff_empty), .Y(dbgpo[23]) );
  OAI21X1 U406 ( .B(n298), .C(n295), .A(n203), .Y(srstz) );
  AND2X1 U407 ( .A(pff_ack[1]), .B(n275), .Y(set04[5]) );
  INVX1 U408 ( .A(n1182), .Y(bus_idle) );
  AND2X1 U409 ( .A(prx_setsta[2]), .B(n14), .Y(set03[2]) );
  AND2X1 U410 ( .A(prx_setsta[1]), .B(n275), .Y(set03[1]) );
  NOR42XL U411 ( .C(n185), .D(n1176), .A(n168), .B(n1149), .Y(n1152) );
  NAND3X1 U412 ( .A(n284), .B(n300), .C(n278), .Y(phyrst) );
  NOR2X1 U413 ( .A(n301), .B(n282), .Y(r_pos_gate) );
  NAND4X1 U414 ( .A(n279), .B(n1176), .C(n1204), .D(n1205), .Y(n1141) );
  NOR2X1 U415 ( .A(n173), .B(n161), .Y(n1204) );
  NOR4XL U416 ( .A(n197), .B(n174), .C(n195), .D(n184), .Y(n1205) );
  NAND3X1 U417 ( .A(n1137), .B(n13), .C(n1134), .Y(upd01) );
  OAI22X1 U418 ( .A(n151), .B(n276), .C(n201), .D(n1127), .Y(wd19[7]) );
  ENOX1 U419 ( .A(n162), .B(n1126), .C(pff_rxpart[0]), .D(n1126), .Y(wd20[0])
         );
  ENOX1 U420 ( .A(n167), .B(n15), .C(pff_rxpart[1]), .D(n1126), .Y(wd20[1]) );
  ENOX1 U421 ( .A(n172), .B(n15), .C(pff_rxpart[2]), .D(n1126), .Y(wd20[2]) );
  ENOX1 U422 ( .A(n179), .B(n15), .C(pff_rxpart[3]), .D(n1126), .Y(wd20[3]) );
  ENOX1 U423 ( .A(n185), .B(n15), .C(pff_rxpart[4]), .D(n1126), .Y(wd20[4]) );
  ENOX1 U424 ( .A(n10), .B(n173), .C(pff_rxpart[10]), .D(n1125), .Y(wd21[2])
         );
  ENOXL U425 ( .A(n1125), .B(n179), .C(pff_rxpart[11]), .D(n1125), .Y(wd21[3])
         );
  ENOX1 U426 ( .A(n10), .B(n184), .C(pff_rxpart[12]), .D(n1125), .Y(wd21[4])
         );
  ENOX1 U427 ( .A(n10), .B(n166), .C(pff_rxpart[9]), .D(n1125), .Y(wd21[1]) );
  ENOX1 U428 ( .A(n10), .B(n190), .C(pff_rxpart[13]), .D(n1125), .Y(wd21[5])
         );
  ENOX1 U429 ( .A(n10), .B(n196), .C(pff_rxpart[14]), .D(n1125), .Y(wd21[6])
         );
  ENOX1 U430 ( .A(n10), .B(n202), .C(pff_rxpart[15]), .D(n1125), .Y(wd21[7])
         );
  ENOX1 U431 ( .A(n161), .B(n1127), .C(inst_ofs_plus[8]), .D(n150), .Y(wd19[0]) );
  ENOX1 U432 ( .A(n167), .B(n1127), .C(inst_ofs_plus[9]), .D(n150), .Y(wd19[1]) );
  ENOX1 U433 ( .A(n172), .B(n1127), .C(inst_ofs_plus[10]), .D(n150), .Y(
        wd19[2]) );
  ENOXL U434 ( .A(n179), .B(n1127), .C(inst_ofs_plus[11]), .D(n150), .Y(
        wd19[3]) );
  ENOX1 U435 ( .A(n185), .B(n1127), .C(inst_ofs_plus[12]), .D(n149), .Y(
        wd19[4]) );
  ENOX1 U436 ( .A(n190), .B(n1127), .C(inst_ofs_plus[13]), .D(n150), .Y(
        wd19[5]) );
  NAND2X1 U437 ( .A(n1139), .B(n15), .Y(upd20) );
  NAND2X1 U438 ( .A(n1139), .B(n10), .Y(upd21) );
  NAND42X1 U439 ( .C(set_hold), .D(cpurst), .A(n1132), .B(n1129), .Y(upd12) );
  AND3X1 U440 ( .A(sfr_r), .B(hit_206), .C(n276), .Y(upd31) );
  AND2X1 U441 ( .A(n266), .B(n273), .Y(hit_206) );
  ENOX1 U442 ( .A(n149), .B(n167), .C(inst_ofs_plus[1]), .D(ictlr_inc), .Y(
        wd18[1]) );
  ENOX1 U443 ( .A(n149), .B(n173), .C(inst_ofs_plus[2]), .D(ictlr_inc), .Y(
        wd18[2]) );
  ENOX1 U444 ( .A(n149), .B(n184), .C(inst_ofs_plus[4]), .D(n150), .Y(wd18[4])
         );
  ENOX1 U445 ( .A(n149), .B(n179), .C(inst_ofs_plus[3]), .D(ictlr_inc), .Y(
        wd18[3]) );
  ENOX1 U446 ( .A(n149), .B(n190), .C(inst_ofs_plus[5]), .D(n150), .Y(wd18[5])
         );
  ENOX1 U447 ( .A(n149), .B(n195), .C(inst_ofs_plus[6]), .D(n150), .Y(wd18[6])
         );
  ENOX1 U448 ( .A(n149), .B(n201), .C(inst_ofs_plus[7]), .D(n150), .Y(wd18[7])
         );
  AND2X1 U449 ( .A(pff_obsd), .B(n275), .Y(set04[3]) );
  NOR2X1 U450 ( .A(n301), .B(n283), .Y(r_osc_lo) );
  AND2X1 U451 ( .A(prx_setsta[4]), .B(n14), .Y(set03[4]) );
  NAND2X1 U452 ( .A(prx_setsta[3]), .B(n275), .Y(n1140) );
  NOR2X1 U453 ( .A(n301), .B(n231), .Y(r_osc_stop) );
  AND2X1 U454 ( .A(i_goidle), .B(n275), .Y(set04[1]) );
  AND2X1 U455 ( .A(i_gobusy), .B(n14), .Y(set04[2]) );
  AND2X1 U456 ( .A(prl_GCTxDone), .B(n14), .Y(set04[6]) );
  AND2X1 U457 ( .A(prl_discard), .B(n275), .Y(set04[7]) );
  XNOR2XL U458 ( .A(n297), .B(N30), .Y(N34) );
  XNOR2XL U459 ( .A(N32), .B(n297), .Y(N33) );
  XOR2X1 U460 ( .A(N30), .B(N29), .Y(N35) );
  XNOR2XL U461 ( .A(N27), .B(N29), .Y(N36) );
  INVX1 U462 ( .A(n1132), .Y(n296) );
  NAND3X1 U463 ( .A(n283), .B(n282), .C(n231), .Y(N81) );
  INVX1 U464 ( .A(n1211), .Y(n294) );
  XNOR2XL U465 ( .A(di_p0[2]), .B(n291), .Y(n1196) );
  XNOR2XL U466 ( .A(di_p0[4]), .B(n289), .Y(n1198) );
  XNOR2XL U467 ( .A(di_p0[6]), .B(n287), .Y(n1200) );
  XNOR2XL U468 ( .A(di_p0[3]), .B(n290), .Y(n1197) );
  XNOR2XL U469 ( .A(di_p0[5]), .B(n288), .Y(n1199) );
  XNOR2XL U470 ( .A(di_p0[7]), .B(n286), .Y(n1201) );
  NAND2X1 U471 ( .A(n203), .B(aswkup), .Y(pwrdn_rstz) );
  BUFX3 U472 ( .A(pff_full), .Y(dbgpo[22]) );
  AND2X1 U473 ( .A(dnchk_en), .B(dm_fault), .Y(dmf_wkup) );
  INVX1 U474 ( .A(n1211), .Y(n1076) );
  MUX2X1 U475 ( .D0(i_pc[2]), .D1(prx_adpn[2]), .S(reg19_7_), .Y(reg30[2]) );
  AND2X1 U476 ( .A(i_pc[6]), .B(n276), .Y(reg30[6]) );
  MUX2X1 U477 ( .D0(s_scp), .D1(m_scp), .S(reg94[5]), .Y(regAD[4]) );
  INVX1 U478 ( .A(n1150), .Y(n238) );
  OAI211X1 U479 ( .C(ictlr_idle), .D(n232), .A(oscdwn_shft[1]), .B(bus_idle), 
        .Y(n1150) );
  AND3X1 U480 ( .A(regD4[1]), .B(n231), .C(n282), .Y(n232) );
  INVX1 U481 ( .A(regD4[0]), .Y(n231) );
  INVX1 U482 ( .A(rstcnt[3]), .Y(n299) );
  INVX1 U483 ( .A(n1189), .Y(n298) );
  OAI211X1 U484 ( .C(rstcnt[2]), .D(rstcnt[1]), .A(n299), .B(rstcnt[4]), .Y(
        n1189) );
  AND3X1 U485 ( .A(hit_207), .B(sfr_r), .C(reg19_7_), .Y(r_psrd) );
  MUX2X1 U486 ( .D0(i_pc[3]), .D1(prx_adpn[3]), .S(reg19_7_), .Y(reg30[3]) );
  MUX2X1 U487 ( .D0(i_pc[0]), .D1(prx_adpn[0]), .S(reg19_7_), .Y(reg30[0]) );
  MUX2X1 U488 ( .D0(i_pc[1]), .D1(prx_adpn[1]), .S(reg19_7_), .Y(reg30[1]) );
  MUX2X1 U489 ( .D0(i_pc[5]), .D1(prx_adpn[5]), .S(reg19_7_), .Y(reg30[5]) );
  MUX2X1 U490 ( .D0(i_pc[4]), .D1(prx_adpn[4]), .S(reg19_7_), .Y(reg30[4]) );
  NAND4X1 U491 ( .A(n1165), .B(n1166), .C(n1167), .D(n1168), .Y(o_intr[1]) );
  AOI22X1 U492 ( .A(reg06[6]), .B(irq04[6]), .C(reg06[7]), .D(irq04[7]), .Y(
        n1165) );
  AOI22X1 U493 ( .A(reg06[0]), .B(irq04[0]), .C(reg06[1]), .D(irq04[1]), .Y(
        n1168) );
  AND2X1 U494 ( .A(i_pc[7]), .B(n276), .Y(reg30[7]) );
  AOI22X1 U495 ( .A(reg06[4]), .B(irq04[4]), .C(reg06[5]), .D(irq04[5]), .Y(
        n1166) );
  OR4X1 U496 ( .A(osc_gate_n[1]), .B(osc_gate_n[0]), .C(osc_gate_n[3]), .D(
        osc_gate_n[2]), .Y(r_osc_gate) );
  INVX1 U497 ( .A(drstz[1]), .Y(n295) );
  MUX2X1 U498 ( .D0(s_ovp), .D1(m_ovp), .S(reg94[4]), .Y(regAD[2]) );
  INVX1 U499 ( .A(reg19_7_), .Y(n276) );
  NAND42X1 U500 ( .C(prl_cany0), .D(n230), .A(i_i2c_idle), .B(n1208), .Y(n1182) );
  INVX1 U501 ( .A(prx_rcvinf[4]), .Y(n230) );
  NOR3XL U502 ( .A(ptx_fsm[0]), .B(ptx_fsm[2]), .C(ptx_fsm[1]), .Y(n1208) );
  NAND4X1 U503 ( .A(n1169), .B(n1170), .C(n1171), .D(n1172), .Y(o_intr[0]) );
  AOI22X1 U504 ( .A(reg05[4]), .B(irq03[4]), .C(reg05[5]), .D(irq03[5]), .Y(
        n1170) );
  AOI22X1 U505 ( .A(reg05[2]), .B(irq03[2]), .C(reg05[3]), .D(irq03[3]), .Y(
        n1171) );
  AOI22X1 U506 ( .A(reg05[6]), .B(irq03[6]), .C(reg05[7]), .D(irq03[7]), .Y(
        n1169) );
  AOI22X1 U507 ( .A(reg05[0]), .B(irq03[0]), .C(reg05[1]), .D(irq03[1]), .Y(
        n1172) );
  INVX1 U508 ( .A(oscdwn_shft[2]), .Y(n301) );
  INVX1 U509 ( .A(regD4[2]), .Y(n282) );
  OAI32X1 U510 ( .A(n1174), .B(i_goidle), .C(n14), .D(r_phyrst[0]), .E(n1175), 
        .Y(n1210) );
  AOI211X1 U511 ( .C(reg11_7_), .D(set03[7]), .A(r_phyrst[1]), .B(n1152), .Y(
        n1175) );
  NAND42X1 U512 ( .C(bkpt_hold), .D(reg12[3]), .A(n231), .B(n282), .Y(
        r_hold_mcu) );
  ENOX1 U513 ( .A(n162), .B(n1123), .C(n1123), .D(lt_reg26_0), .Y(
        i2c_mode_wdat) );
  AOI21X1 U514 ( .B(n1181), .C(n1123), .A(n1182), .Y(i2c_mode_upd) );
  XNOR2XL U515 ( .A(r_hwi2c_en), .B(lt_reg26_0), .Y(n1181) );
  OAI21X1 U516 ( .B(r_fifopop), .C(r_fifopsh), .A(r_first), .Y(n1137) );
  OAI21BBX1 U517 ( .A(n296), .B(reg12[3]), .C(n1131), .Y(wd12[3]) );
  AOI32XL U518 ( .A(n1132), .B(n1129), .C(set_hold), .D(n1133), .E(n174), .Y(
        n1131) );
  NOR21XL U519 ( .B(n1137), .A(n1138), .Y(wd01[6]) );
  AOI22X1 U520 ( .A(r_first), .B(n1136), .C(n280), .D(n194), .Y(n1138) );
  NOR21XL U521 ( .B(n1134), .A(n1135), .Y(wd01[7]) );
  AOI22X1 U522 ( .A(r_last), .B(n1136), .C(n280), .D(n200), .Y(n1135) );
  OAI21X1 U523 ( .B(n185), .C(n1129), .A(n1130), .Y(wd12[4]) );
  AOI21X1 U524 ( .B(reg12[4]), .C(n1129), .A(n296), .Y(n1130) );
  OAI21X1 U525 ( .B(n1203), .C(n1182), .A(n1141), .Y(N23) );
  NOR21XL U526 ( .B(n1142), .A(rstcnt[4]), .Y(n1203) );
  ENOX1 U527 ( .A(n190), .B(n15), .C(pff_rxpart[5]), .D(n1126), .Y(wd20[5]) );
  ENOX1 U528 ( .A(n196), .B(n15), .C(pff_rxpart[6]), .D(n1126), .Y(wd20[6]) );
  ENOX1 U529 ( .A(n202), .B(n15), .C(pff_rxpart[7]), .D(n1126), .Y(wd20[7]) );
  AO22AXL U530 ( .A(r_pshords), .B(n281), .C(sfr_wdat[0]), .D(n281), .Y(
        wd12[0]) );
  ENOX1 U531 ( .A(n167), .B(n281), .C(reg12_1), .D(n281), .Y(wd12[1]) );
  AO22AXL U532 ( .A(r_txshrt), .B(n281), .C(sfr_wdat[2]), .D(n281), .Y(wd12[2]) );
  ENOX1 U533 ( .A(n190), .B(n281), .C(reg12[5]), .D(n281), .Y(wd12[5]) );
  ENOX1 U534 ( .A(n195), .B(n11), .C(reg12[6]), .D(n281), .Y(wd12[6]) );
  ENOX1 U535 ( .A(n202), .B(n11), .C(reg12[7]), .D(n281), .Y(wd12[7]) );
  ENOX1 U536 ( .A(n10), .B(n162), .C(pff_rxpart[8]), .D(n1125), .Y(wd21[0]) );
  ENOX1 U537 ( .A(n196), .B(n1127), .C(inst_ofs_plus[14]), .D(n150), .Y(
        wd19[6]) );
  ENOX1 U538 ( .A(n185), .B(n13), .C(r_txnumk[4]), .D(n1136), .Y(wd01[4]) );
  ENOX1 U539 ( .A(n190), .B(n13), .C(r_unlock), .D(n1136), .Y(wd01[5]) );
  NAND2X1 U540 ( .A(r_last), .B(r_fifopsh), .Y(n1134) );
  NAND3X1 U541 ( .A(n1178), .B(n1179), .C(n1180), .Y(i2c_stretch) );
  AOI22X1 U542 ( .A(reg28[2]), .B(reg27[2]), .C(reg28[3]), .D(reg27[3]), .Y(
        n1178) );
  AOI22X1 U543 ( .A(reg28[0]), .B(reg27[0]), .C(reg28[1]), .D(reg27[1]), .Y(
        n1179) );
  AOI222XL U544 ( .A(reg28[7]), .B(reg27[7]), .C(reg28[4]), .D(reg27[4]), .E(
        reg28[6]), .F(reg27[6]), .Y(n1180) );
  ENOX1 U545 ( .A(n149), .B(n161), .C(inst_ofs_plus[0]), .D(n149), .Y(wd18[0])
         );
  AOI22X1 U546 ( .A(reg06[2]), .B(irq04[2]), .C(reg06[3]), .D(irq04[3]), .Y(
        n1167) );
  INVX1 U547 ( .A(regD4[1]), .Y(n283) );
  NOR21XL U548 ( .B(prx_setsta[6]), .A(prl_cany0), .Y(set03[6]) );
  AOI21BBXL U549 ( .B(r_auto_gdcrc[1]), .C(n1140), .A(set03[6]), .Y(n1139) );
  AO21X1 U550 ( .B(n1144), .C(n1145), .A(reg11_4), .Y(r_rxords_ena[4]) );
  NOR3XL U551 ( .A(r_rxords_ena[0]), .B(r_rxords_ena[2]), .C(r_rxords_ena[1]), 
        .Y(n1144) );
  NOR3XL U552 ( .A(r_rxords_ena[3]), .B(r_rxords_ena[6]), .C(r_rxords_ena[5]), 
        .Y(n1145) );
  OAI31XL U553 ( .A(n295), .B(r_phyrst[1]), .C(n298), .D(n203), .Y(prstz) );
  AND2X1 U554 ( .A(prx_setsta[5]), .B(n275), .Y(set03[5]) );
  AOI22X1 U555 ( .A(reg27[6]), .B(irq28[6]), .C(reg27[7]), .D(irq28[7]), .Y(
        n1161) );
  NAND4X1 U556 ( .A(n1161), .B(n1162), .C(n1163), .D(n1164), .Y(o_intr[2]) );
  AOI22X1 U557 ( .A(reg27[4]), .B(irq28[4]), .C(reg27[5]), .D(irq28[5]), .Y(
        n1162) );
  AOI22X1 U558 ( .A(reg27[0]), .B(irq28[0]), .C(reg27[1]), .D(irq28[1]), .Y(
        n1164) );
  NOR21XL U559 ( .B(regD4[4]), .A(n301), .Y(r_ocdrv_enz) );
  AND2X1 U560 ( .A(ptx_ack), .B(n275), .Y(set04[0]) );
  AOI22X1 U561 ( .A(reg27[2]), .B(irq28[2]), .C(reg27[3]), .D(irq28[3]), .Y(
        n1163) );
  AOI221XL U562 ( .A(regAF[2]), .B(regAE[2]), .C(regAF[4]), .D(regAE[4]), .E(
        n285), .Y(r_srcctl[0]) );
  INVX1 U563 ( .A(regE3_0), .Y(n285) );
  AND2X1 U564 ( .A(reg94[7]), .B(reg94[6]), .Y(r_otpi_gate) );
  AO22AXL U565 ( .A(reg94[4]), .B(m_ovp_sta), .C(s_ovp_sta), .D(reg94[4]), .Y(
        setAE[2]) );
  AO22AXL U566 ( .A(reg94[5]), .B(m_scp_sta), .C(s_scp_sta), .D(reg94[5]), .Y(
        setAE[4]) );
  NOR21XL U567 ( .B(regD4[3]), .A(n301), .Y(r_pwrdn) );
  NAND4X1 U568 ( .A(n1153), .B(n1154), .C(n1155), .D(n1156), .Y(o_intr[4]) );
  AOI22X1 U569 ( .A(regAF[6]), .B(irqAE[6]), .C(regAF[7]), .D(irqAE[7]), .Y(
        n1153) );
  AOI22X1 U570 ( .A(regAF[0]), .B(irqAE[0]), .C(regAF[1]), .D(irqAE[1]), .Y(
        n1156) );
  AOI22X1 U571 ( .A(irqAE[2]), .B(regAF[2]), .C(regAF[3]), .D(irqAE[3]), .Y(
        n1155) );
  AOI22X1 U572 ( .A(irqAE[4]), .B(regAF[4]), .C(irqAE[5]), .D(regAF[5]), .Y(
        n1154) );
  XNOR2XL U573 ( .A(d_p0[0]), .B(n293), .Y(setDF[0]) );
  XNOR2XL U574 ( .A(d_p0[1]), .B(n292), .Y(setDF[1]) );
  XNOR2XL U575 ( .A(d_p0[2]), .B(n291), .Y(setDF[2]) );
  XNOR2XL U576 ( .A(d_p0[3]), .B(n290), .Y(setDF[3]) );
  XNOR2XL U577 ( .A(d_p0[4]), .B(n289), .Y(setDF[4]) );
  INVX1 U578 ( .A(prl_cany0), .Y(n275) );
  XNOR2XL U579 ( .A(rstcnt[4]), .B(n299), .Y(N24) );
  XNOR2XL U580 ( .A(n1202), .B(N24), .Y(N26) );
  XNOR2XL U581 ( .A(rstcnt[2]), .B(rstcnt[1]), .Y(n1202) );
  AND2X1 U582 ( .A(prx_setsta[0]), .B(n275), .Y(set03[0]) );
  XOR2X1 U583 ( .A(N26), .B(rstcnt[0]), .Y(N27) );
  XOR2X1 U584 ( .A(rstcnt[2]), .B(N24), .Y(N25) );
  NOR42XL U585 ( .C(n1206), .D(r_inst_ofs[10]), .A(r_inst_ofs[8]), .B(n1207), 
        .Y(n1176) );
  NAND4X1 U586 ( .A(r_inst_ofs[14]), .B(r_inst_ofs[13]), .C(r_inst_ofs[12]), 
        .D(r_inst_ofs[11]), .Y(n1207) );
  NOR2X1 U587 ( .A(reg19_7_), .B(r_inst_ofs[9]), .Y(n1206) );
  AOI22X1 U588 ( .A(regDE[0]), .B(irqDF[0]), .C(regDE[1]), .D(irqDF[1]), .Y(
        n1160) );
  AOI22X1 U589 ( .A(regDE[2]), .B(irqDF[2]), .C(regDE[3]), .D(irqDF[3]), .Y(
        n1159) );
  XNOR2XL U590 ( .A(d_p0[6]), .B(n287), .Y(setDF[6]) );
  XNOR2XL U591 ( .A(d_p0[7]), .B(n286), .Y(setDF[7]) );
  XNOR2XL U592 ( .A(d_p0[5]), .B(n288), .Y(setDF[5]) );
  NAND4X1 U593 ( .A(n1157), .B(n1158), .C(n1159), .D(n1160), .Y(o_intr[3]) );
  AOI22X1 U594 ( .A(regDE[6]), .B(irqDF[6]), .C(regDE[7]), .D(irqDF[7]), .Y(
        n1157) );
  AOI22X1 U595 ( .A(regDE[4]), .B(irqDF[4]), .C(regDE[5]), .D(irqDF[5]), .Y(
        n1158) );
  INVX1 U596 ( .A(ff_p0[2]), .Y(n291) );
  INVX1 U597 ( .A(ff_p0[6]), .Y(n287) );
  INVX1 U598 ( .A(ff_p0[5]), .Y(n288) );
  INVX1 U599 ( .A(ff_p0[7]), .Y(n286) );
  INVX1 U600 ( .A(ff_p0[0]), .Y(n293) );
  INVX1 U601 ( .A(ff_p0[1]), .Y(n292) );
  INVX1 U602 ( .A(ff_p0[3]), .Y(n290) );
  INVX1 U603 ( .A(ff_p0[4]), .Y(n289) );
  OAI22X1 U604 ( .A(r_phyrst[0]), .B(n300), .C(n1173), .D(n1174), .Y(n1209) );
  NOR2X1 U605 ( .A(i_goidle), .B(n14), .Y(n1173) );
  INVX1 U606 ( .A(reg25_0_), .Y(r_i2c_ninc) );
  NAND2X1 U607 ( .A(rstcnt[4]), .B(n1142), .Y(n1132) );
  NOR4XL U608 ( .A(rstcnt[0]), .B(rstcnt[1]), .C(rstcnt[2]), .D(rstcnt[3]), 
        .Y(n1142) );
  INVX1 U609 ( .A(r_phyrst[1]), .Y(n300) );
  NAND2X1 U610 ( .A(r_phyrst[0]), .B(n300), .Y(n1174) );
  NAND42X1 U611 ( .C(di_stbovp_clr), .D(di_rd_det_clr), .A(n294), .B(n1188), 
        .Y(aswkup) );
  NOR3XL U612 ( .A(dm_fault_clr), .B(p0_chg_clr), .C(i_tmrf), .Y(n1188) );
  AND2X1 U613 ( .A(regE3[3]), .B(n1143), .Y(r_srcctl[3]) );
  AND2X1 U614 ( .A(regE3[2]), .B(n1143), .Y(r_srcctl[2]) );
  INVX1 U615 ( .A(regD3_3), .Y(r_gpio_ie[0]) );
  NAND2X1 U616 ( .A(srstz), .B(n7), .Y(n1211) );
  OAI21X1 U617 ( .B(osc_low_clr), .C(n1211), .A(n203), .Y(osc_low_rstz) );
  AOI22X1 U618 ( .A(regDE[0]), .B(n1194), .C(regDE[1]), .D(n1195), .Y(n1193)
         );
  XNOR2XL U619 ( .A(di_p0[1]), .B(n292), .Y(n1195) );
  XNOR2XL U620 ( .A(di_p0[0]), .B(n293), .Y(n1194) );
  AOI22X1 U621 ( .A(regAF[5]), .B(regAE[5]), .C(regAD[5]), .D(i_vcbyval), .Y(
        n1143) );
  INVX1 U622 ( .A(regD3_7_), .Y(r_gpio_ie[1]) );
  NAND4X1 U623 ( .A(n1190), .B(n1191), .C(n1192), .D(n1193), .Y(as_p0_chg) );
  AOI22X1 U624 ( .A(regDE[6]), .B(n1200), .C(regDE[7]), .D(n1201), .Y(n1190)
         );
  AOI22X1 U625 ( .A(regDE[4]), .B(n1198), .C(regDE[5]), .D(n1199), .Y(n1191)
         );
  AOI22X1 U626 ( .A(regDE[2]), .B(n1196), .C(regDE[3]), .D(n1197), .Y(n1192)
         );
  INVX1 U627 ( .A(sfr_addr[7]), .Y(n206) );
  BUFX3 U628 ( .A(sfr_w), .Y(n71) );
  BUFXL U629 ( .A(sfr_w), .Y(n72) );
  NAND21X1 U630 ( .B(n154), .A(n31), .Y(n234) );
  NAND32XL U631 ( .B(n255), .C(n154), .A(n156), .Y(n256) );
  NAND32XL U632 ( .B(n241), .C(n154), .A(n156), .Y(n211) );
  NAND32XL U633 ( .B(n154), .C(n155), .A(n209), .Y(n210) );
  NAND21X1 U634 ( .B(n154), .A(n62), .Y(n208) );
  NAND43X1 U635 ( .B(n153), .C(n242), .D(n156), .A(n241), .Y(n243) );
  NAND43X1 U636 ( .B(n153), .C(n155), .D(n242), .A(n236), .Y(n237) );
  NOR2X1 U637 ( .A(n155), .B(n153), .Y(n302) );
  INVXL U638 ( .A(sfr_addr[5]), .Y(n154) );
  OAI21BBXL U639 ( .A(hit_194), .B(n72), .C(n151), .Y(upd18) );
  NOR32XL U640 ( .B(hit_207), .C(n71), .A(n276), .Y(r_pswr) );
  AND3X2 U641 ( .A(n274), .B(n174), .C(n238), .Y(ps_pwrdn) );
  NAND21XL U642 ( .B(n258), .A(n259), .Y(n1126) );
  NAND21XL U643 ( .B(n258), .A(n265), .Y(n1129) );
  NAND21XL U644 ( .B(n258), .A(n266), .Y(n1185) );
  NAND21XL U645 ( .B(n258), .A(n264), .Y(n1186) );
  AND4XL U646 ( .A(n215), .B(n155), .C(n263), .D(n153), .Y(we_232) );
  NAND21XL U647 ( .B(n153), .A(n62), .Y(n257) );
  NAND32XL U648 ( .B(n157), .C(n255), .A(n153), .Y(n233) );
  NAND21XL U649 ( .B(n153), .A(n31), .Y(n217) );
  XOR2X1 U650 ( .A(add_179_carry[4]), .B(rstcnt[4]), .Y(N32) );
endmodule


module regbank_a0_DW_rightsh_0 ( A, DATA_TC, SH, B );
  input [1023:0] A;
  input [9:0] SH;
  output [1023:0] B;
  input DATA_TC;
  wire   n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611,
         n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621,
         n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631,
         n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641,
         n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651,
         n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661,
         n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671,
         n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681,
         n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691,
         n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701,
         n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711,
         n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721,
         n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731,
         n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741,
         n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751,
         n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761,
         n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771,
         n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781,
         n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791,
         n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801,
         n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811,
         n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821,
         n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831,
         n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841,
         n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851,
         n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861,
         n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871,
         n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881,
         n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891,
         n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901,
         n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911,
         n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921,
         n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931,
         n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941,
         n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951,
         n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961,
         n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971,
         n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981,
         n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991,
         n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001,
         n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011,
         n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021,
         n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031,
         n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041,
         n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051,
         n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061,
         n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071,
         n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081,
         n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091,
         n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101,
         n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111,
         n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121,
         n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131,
         n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141,
         n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151,
         n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161,
         n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171,
         n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181,
         n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191,
         n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201,
         n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211,
         n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221,
         n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231,
         n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241,
         n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251,
         n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261,
         n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271,
         n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281,
         n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291,
         n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301,
         n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311,
         n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321,
         n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329;

  BUFX3 U2565 ( .A(n3757), .Y(n3602) );
  INVXL U2566 ( .A(n3768), .Y(n3757) );
  INVX1 U2567 ( .A(n3629), .Y(n3653) );
  MUX2IXL U2568 ( .D0(n4305), .D1(n4306), .S(n3611), .Y(n4304) );
  NAND2XL U2569 ( .A(n4213), .B(n3611), .Y(n4209) );
  MUX2IXL U2570 ( .D0(n4263), .D1(n4264), .S(n3607), .Y(n4262) );
  MUX2IXL U2571 ( .D0(n3929), .D1(n3930), .S(n3607), .Y(n3928) );
  MUX4XL U2572 ( .D0(n3900), .D1(n3901), .D2(n3902), .D3(n3903), .S0(n3607), 
        .S1(n3664), .Y(n3899) );
  MUX2IXL U2573 ( .D0(n4002), .D1(n4003), .S(n3607), .Y(n4001) );
  MUX2IXL U2574 ( .D0(n4009), .D1(n4010), .S(n3607), .Y(n4008) );
  INVX20 U2575 ( .A(n3635), .Y(n3767) );
  INVX2 U2576 ( .A(SH[9]), .Y(n3635) );
  INVX20 U2577 ( .A(n3635), .Y(n3756) );
  BUFX3 U2578 ( .A(n3754), .Y(n3603) );
  INVXL U2579 ( .A(n3635), .Y(n3754) );
  INVX20 U2580 ( .A(n3635), .Y(n3753) );
  INVX3 U2581 ( .A(n3605), .Y(n3606) );
  INVX2 U2582 ( .A(n3605), .Y(n3607) );
  BUFX6 U2583 ( .A(n3761), .Y(n3604) );
  INVX2 U2584 ( .A(n3755), .Y(n3605) );
  INVX1 U2585 ( .A(n3706), .Y(n3690) );
  INVX1 U2586 ( .A(n3709), .Y(n3693) );
  MUX2X1 U2587 ( .D0(n4199), .D1(n4200), .S(n3673), .Y(n3622) );
  MUX2X1 U2588 ( .D0(n4221), .D1(n4220), .S(n3676), .Y(n3621) );
  MUX2X1 U2589 ( .D0(n3984), .D1(n3985), .S(SH[7]), .Y(B[4]) );
  MUX2X1 U2590 ( .D0(n3947), .D1(n3948), .S(n3681), .Y(n3628) );
  MUX2X1 U2591 ( .D0(n4285), .D1(n4286), .S(n3672), .Y(n3633) );
  MUX2X1 U2592 ( .D0(n3613), .D1(n3614), .S(n3673), .Y(n3630) );
  INVX2 U2593 ( .A(SH[5]), .Y(n3680) );
  INVX1 U2594 ( .A(SH[8]), .Y(n3751) );
  INVX1 U2595 ( .A(SH[9]), .Y(n3768) );
  MUX2X1 U2596 ( .D0(n3608), .D1(n3609), .S(SH[7]), .Y(B[3]) );
  MUX2IX1 U2597 ( .D0(n4088), .D1(n4089), .S(n3681), .Y(n3608) );
  MUX4X1 U2598 ( .D0(n4057), .D1(n4058), .D2(n4059), .D3(n4060), .S0(n3678), 
        .S1(n3682), .Y(n3609) );
  INVXL U2599 ( .A(n3629), .Y(n3762) );
  INVXL U2600 ( .A(n3768), .Y(n3763) );
  INVX1 U2601 ( .A(n3709), .Y(n3689) );
  INVXL U2602 ( .A(n3635), .Y(n3610) );
  INVX1 U2603 ( .A(n3710), .Y(n3688) );
  INVX1 U2604 ( .A(n3670), .Y(n3658) );
  INVX1 U2605 ( .A(n3635), .Y(n3611) );
  INVXL U2606 ( .A(n3710), .Y(n3687) );
  INVX1 U2607 ( .A(n3670), .Y(n3659) );
  MUX4XL U2608 ( .D0(A[241]), .D1(A[753]), .D2(A[497]), .D3(A[1009]), .S0(
        n3648), .S1(n3699), .Y(n4201) );
  MUX4XL U2609 ( .D0(n4094), .D1(n4095), .D2(n4096), .D3(n4097), .S0(n3658), 
        .S1(n3602), .Y(n4093) );
  MUX4XL U2610 ( .D0(n4203), .D1(n4204), .D2(n4205), .D3(n4206), .S0(n3658), 
        .S1(n3602), .Y(n4199) );
  MUX4XL U2611 ( .D0(n4299), .D1(n4300), .D2(n4301), .D3(n4302), .S0(n3658), 
        .S1(n3766), .Y(n4298) );
  MUX4XL U2612 ( .D0(n3811), .D1(n3812), .D2(n3813), .D3(n3814), .S0(n3658), 
        .S1(n3606), .Y(n3810) );
  INVX1 U2613 ( .A(n3709), .Y(n3691) );
  INVX1 U2614 ( .A(n3676), .Y(n3671) );
  INVX1 U2615 ( .A(n3629), .Y(n3760) );
  INVX1 U2616 ( .A(n3668), .Y(n3666) );
  INVXL U2617 ( .A(n3668), .Y(n3667) );
  INVXL U2618 ( .A(n3708), .Y(n3695) );
  INVXL U2619 ( .A(n3676), .Y(n3672) );
  INVXL U2620 ( .A(n3708), .Y(n3694) );
  INVXL U2621 ( .A(n3668), .Y(n3665) );
  INVXL U2622 ( .A(n3708), .Y(n3696) );
  INVX1 U2623 ( .A(n3676), .Y(n3674) );
  INVX3 U2624 ( .A(n3711), .Y(n3685) );
  INVXL U2625 ( .A(n3668), .Y(n3664) );
  INVXL U2626 ( .A(n3668), .Y(n3663) );
  INVX1 U2627 ( .A(n3750), .Y(n3707) );
  INVX1 U2628 ( .A(n3683), .Y(n3682) );
  INVX1 U2629 ( .A(n3683), .Y(n3681) );
  INVXL U2630 ( .A(n3676), .Y(n3673) );
  INVXL U2631 ( .A(SH[8]), .Y(n3625) );
  MUX2IXL U2632 ( .D0(n4071), .D1(n4072), .S(n3653), .Y(n3615) );
  MUX2IX1 U2633 ( .D0(n4266), .D1(n4267), .S(n3660), .Y(n3614) );
  MUX2IX1 U2634 ( .D0(A[223]), .D1(A[479]), .S(n3691), .Y(n3787) );
  NAND21XL U2635 ( .B(n3619), .A(n3603), .Y(n4070) );
  MUX2XL U2636 ( .D0(A[715]), .D1(A[971]), .S(n3747), .Y(n3619) );
  INVXL U2637 ( .A(n3635), .Y(n3755) );
  INVXL U2638 ( .A(n3768), .Y(n3766) );
  INVXL U2639 ( .A(n3635), .Y(n3761) );
  INVXL U2640 ( .A(n3768), .Y(n3648) );
  INVXL U2641 ( .A(n3676), .Y(n3675) );
  MUX2IX1 U2642 ( .D0(n3612), .D1(n4061), .S(n3673), .Y(n4060) );
  MUX4XL U2643 ( .D0(n4064), .D1(n4065), .D2(n4066), .D3(n4067), .S0(n3658), 
        .S1(n3606), .Y(n3612) );
  MUX4XL U2644 ( .D0(n4268), .D1(n4269), .D2(n4270), .D3(n4271), .S0(n3658), 
        .S1(n3753), .Y(n3613) );
  MUX4X1 U2645 ( .D0(n4068), .D1(n4069), .D2(n4070), .D3(n3615), .S0(n3672), 
        .S1(n3663), .Y(n4059) );
  MUX4X1 U2646 ( .D0(n3630), .D1(n3631), .D2(n3632), .D3(n3633), .S0(n3680), 
        .S1(n3683), .Y(n3617) );
  MUX2BX1 U2647 ( .D0(n4265), .D1(n3617), .S(SH[7]), .Y(B[0]) );
  INVXL U2648 ( .A(A[500]), .Y(n3651) );
  MUX4XL U2649 ( .D0(A[254]), .D1(A[766]), .D2(A[510]), .D3(A[1022]), .S0(
        n3624), .S1(n3700), .Y(n3851) );
  MUX2IXL U2650 ( .D0(A[221]), .D1(A[477]), .S(n3694), .Y(n3929) );
  MUX2XL U2651 ( .D0(A[128]), .D1(A[384]), .S(n3684), .Y(n3616) );
  MUX2IXL U2652 ( .D0(A[717]), .D1(A[973]), .S(n3693), .Y(n3931) );
  MUX2IXL U2653 ( .D0(A[222]), .D1(A[478]), .S(n3692), .Y(n3860) );
  MUX2IXL U2654 ( .D0(A[714]), .D1(A[970]), .S(n3687), .Y(n4145) );
  NOR2XL U2655 ( .A(A[287]), .B(n3734), .Y(n3835) );
  NOR2XL U2656 ( .A(A[286]), .B(n3734), .Y(n3906) );
  NOR2XL U2657 ( .A(A[310]), .B(n3734), .Y(n3900) );
  MUX2IXL U2658 ( .D0(A[718]), .D1(A[974]), .S(n3692), .Y(n3862) );
  INVX1 U2659 ( .A(n3629), .Y(n3758) );
  INVX1 U2660 ( .A(SH[9]), .Y(n3629) );
  INVX1 U2661 ( .A(n3604), .Y(n3764) );
  INVX1 U2662 ( .A(n3648), .Y(n3765) );
  INVX1 U2663 ( .A(n3709), .Y(n3692) );
  INVX3 U2664 ( .A(n3711), .Y(n3684) );
  INVX1 U2665 ( .A(n3635), .Y(n3759) );
  INVX1 U2666 ( .A(n3680), .Y(n3678) );
  INVX1 U2667 ( .A(n3707), .Y(n3699) );
  INVX1 U2668 ( .A(n3680), .Y(n3677) );
  INVX1 U2669 ( .A(n3707), .Y(n3697) );
  INVX1 U2670 ( .A(n3669), .Y(n3661) );
  INVX1 U2671 ( .A(n3707), .Y(n3698) );
  INVX1 U2672 ( .A(n3669), .Y(n3660) );
  INVX1 U2673 ( .A(n3669), .Y(n3662) );
  INVXL U2674 ( .A(n3705), .Y(n3701) );
  INVXL U2675 ( .A(n3705), .Y(n3702) );
  INVX1 U2676 ( .A(n3680), .Y(n3679) );
  INVX1 U2677 ( .A(n3625), .Y(n3742) );
  INVX1 U2678 ( .A(n3625), .Y(n3747) );
  INVX1 U2679 ( .A(n3625), .Y(n3746) );
  INVX1 U2680 ( .A(n3625), .Y(n3743) );
  INVX1 U2681 ( .A(SH[3]), .Y(n3668) );
  INVX1 U2682 ( .A(SH[3]), .Y(n3669) );
  INVX1 U2683 ( .A(SH[3]), .Y(n3670) );
  INVX1 U2684 ( .A(n3625), .Y(n3744) );
  INVX1 U2685 ( .A(SH[6]), .Y(n3683) );
  INVX1 U2686 ( .A(SH[4]), .Y(n3676) );
  INVX1 U2687 ( .A(A[1012]), .Y(n3652) );
  INVX1 U2688 ( .A(A[1020]), .Y(n3647) );
  NAND21XL U2689 ( .B(n3616), .A(n3764), .Y(n4291) );
  MUX2BX1 U2690 ( .D0(n4198), .D1(n3618), .S(SH[7]), .Y(B[1]) );
  MUX4X1 U2691 ( .D0(n3620), .D1(n3621), .D2(n3622), .D3(n3623), .S0(n3680), 
        .S1(n3682), .Y(n3618) );
  MUX2IX1 U2692 ( .D0(n3628), .D1(n3627), .S(SH[7]), .Y(B[5]) );
  INVX1 U2693 ( .A(A[932]), .Y(n3643) );
  INVX1 U2694 ( .A(A[676]), .Y(n3641) );
  INVX1 U2695 ( .A(A[420]), .Y(n3642) );
  INVX1 U2696 ( .A(A[244]), .Y(n3649) );
  INVX1 U2697 ( .A(A[756]), .Y(n3650) );
  INVX1 U2698 ( .A(A[929]), .Y(n3657) );
  INVX1 U2699 ( .A(A[508]), .Y(n3646) );
  INVX1 U2700 ( .A(A[161]), .Y(n3654) );
  INVX1 U2701 ( .A(A[764]), .Y(n3645) );
  INVX1 U2702 ( .A(A[252]), .Y(n3644) );
  INVX1 U2703 ( .A(A[417]), .Y(n3656) );
  INVX1 U2704 ( .A(A[164]), .Y(n3640) );
  INVX1 U2705 ( .A(A[673]), .Y(n3655) );
  INVX1 U2706 ( .A(A[940]), .Y(n3639) );
  INVX1 U2707 ( .A(A[172]), .Y(n3636) );
  INVX1 U2708 ( .A(A[684]), .Y(n3637) );
  INVX1 U2709 ( .A(A[428]), .Y(n3638) );
  MUX4X1 U2710 ( .D0(A[179]), .D1(A[691]), .D2(A[435]), .D3(A[947]), .S0(n3756), .S1(n3696), .Y(n4074) );
  MUX4IX1 U2711 ( .D0(n4214), .D1(n4215), .D2(n4216), .D3(n4217), .S0(n3671), 
        .S1(n3665), .Y(n3620) );
  MUX4IX1 U2712 ( .D0(n4207), .D1(n4208), .D2(n4209), .D3(n4210), .S0(n3672), 
        .S1(n3666), .Y(n3623) );
  INVXL U2713 ( .A(n3768), .Y(n3624) );
  MUX4IX1 U2714 ( .D0(n3656), .D1(n3657), .D2(n3654), .D3(n3655), .S0(n3766), 
        .S1(n3625), .Y(n4214) );
  NOR2XL U2715 ( .A(A[1007]), .B(n3711), .Y(n3782) );
  INVX1 U2716 ( .A(n3706), .Y(n3700) );
  INVX2 U2717 ( .A(n3710), .Y(n3686) );
  INVX1 U2718 ( .A(n3706), .Y(n3704) );
  INVX1 U2719 ( .A(n3711), .Y(n3703) );
  MUX4XL U2720 ( .D0(A[137]), .D1(A[649]), .D2(A[393]), .D3(A[905]), .S0(n3610), .S1(n3745), .Y(n3626) );
  MUX2IX1 U2721 ( .D0(n3626), .D1(n4226), .S(n3669), .Y(n4220) );
  MUX2IXL U2722 ( .D0(n4161), .D1(n4162), .S(n3681), .Y(n4125) );
  MUX4IX1 U2723 ( .D0(n3913), .D1(n3914), .D2(n3915), .D3(n3916), .S0(n3677), 
        .S1(n3681), .Y(n3627) );
  MUX4XL U2724 ( .D0(n3863), .D1(n3864), .D2(n3865), .D3(n3866), .S0(n3671), 
        .S1(n3665), .Y(n3845) );
  MUX2IXL U2725 ( .D0(n3867), .D1(n3868), .S(n3756), .Y(n3866) );
  MUX4IXL U2726 ( .D0(n4272), .D1(n4273), .D2(n4274), .D3(n4275), .S0(n3672), 
        .S1(n3666), .Y(n3631) );
  MUX4IX1 U2727 ( .D0(n4279), .D1(n4280), .D2(n4281), .D3(n4282), .S0(n3671), 
        .S1(n3667), .Y(n3632) );
  INVXL U2728 ( .A(n3606), .Y(n3634) );
  INVX1 U2729 ( .A(n3625), .Y(n3740) );
  INVX1 U2730 ( .A(n3625), .Y(n3748) );
  INVX1 U2731 ( .A(n3625), .Y(n3741) );
  INVX1 U2732 ( .A(n3625), .Y(n3745) );
  INVX1 U2733 ( .A(n3752), .Y(n3750) );
  INVX1 U2734 ( .A(n3751), .Y(n3749) );
  INVXL U2735 ( .A(n3740), .Y(n3739) );
  INVXL U2736 ( .A(n3748), .Y(n3714) );
  INVXL U2737 ( .A(n3748), .Y(n3713) );
  INVXL U2738 ( .A(n3748), .Y(n3712) );
  INVXL U2739 ( .A(n3747), .Y(n3717) );
  INVX1 U2740 ( .A(n3747), .Y(n3716) );
  INVX1 U2741 ( .A(n3747), .Y(n3715) );
  INVX1 U2742 ( .A(n3746), .Y(n3720) );
  INVX1 U2743 ( .A(n3746), .Y(n3719) );
  INVXL U2744 ( .A(n3746), .Y(n3718) );
  INVXL U2745 ( .A(n3743), .Y(n3732) );
  INVX1 U2746 ( .A(n3743), .Y(n3731) );
  INVX1 U2747 ( .A(n3743), .Y(n3730) );
  INVX1 U2748 ( .A(n3742), .Y(n3735) );
  INVX1 U2749 ( .A(n3742), .Y(n3734) );
  INVX1 U2750 ( .A(n3742), .Y(n3733) );
  INVX1 U2751 ( .A(n3741), .Y(n3738) );
  INVX1 U2752 ( .A(n3741), .Y(n3737) );
  INVXL U2753 ( .A(n3741), .Y(n3736) );
  INVXL U2754 ( .A(n3745), .Y(n3723) );
  INVXL U2755 ( .A(n3745), .Y(n3722) );
  INVXL U2756 ( .A(n3745), .Y(n3721) );
  INVXL U2757 ( .A(n3744), .Y(n3726) );
  INVXL U2758 ( .A(n3744), .Y(n3725) );
  INVXL U2759 ( .A(n3744), .Y(n3724) );
  INVXL U2760 ( .A(n3704), .Y(n3729) );
  INVXL U2761 ( .A(n3704), .Y(n3728) );
  INVXL U2762 ( .A(n3750), .Y(n3727) );
  INVX1 U2763 ( .A(SH[8]), .Y(n3706) );
  INVX1 U2764 ( .A(n3750), .Y(n3705) );
  INVX1 U2765 ( .A(n3749), .Y(n3709) );
  INVXL U2766 ( .A(n3749), .Y(n3711) );
  INVX1 U2767 ( .A(SH[8]), .Y(n3710) );
  MUX2IX1 U2768 ( .D0(n4202), .D1(n4201), .S(n3669), .Y(n4200) );
  MUX4IXL U2769 ( .D0(n3637), .D1(n3636), .D2(n3639), .D3(n3638), .S0(n3629), 
        .S1(n3694), .Y(n4007) );
  MUX4X1 U2770 ( .D0(A[181]), .D1(A[693]), .D2(A[437]), .D3(A[949]), .S0(n3754), .S1(n3696), .Y(n3933) );
  MUX4IX1 U2771 ( .D0(n3640), .D1(n3641), .D2(n3642), .D3(n3643), .S0(n3753), 
        .S1(n3694), .Y(n4005) );
  MUX4IX1 U2772 ( .D0(n3644), .D1(n3645), .D2(n3646), .D3(n3647), .S0(n3611), 
        .S1(n3699), .Y(n3993) );
  MUX4IX1 U2773 ( .D0(n3649), .D1(n3650), .D2(n3651), .D3(n3652), .S0(n3760), 
        .S1(n3698), .Y(n3992) );
  MUX2IX1 U2774 ( .D0(n3993), .D1(n3992), .S(n3669), .Y(n3991) );
  INVXL U2775 ( .A(SH[8]), .Y(n3752) );
  NAND31XL U2776 ( .C(A[981]), .A(n3742), .B(n3762), .Y(n3926) );
  MUX4XL U2777 ( .D0(n4175), .D1(n4176), .D2(n4177), .D3(n4178), .S0(n3653), 
        .S1(n3665), .Y(n4164) );
  MUX4XL U2778 ( .D0(n4154), .D1(n4155), .D2(n4156), .D3(n4157), .S0(n3653), 
        .S1(n3665), .Y(n4153) );
  MUX4XL U2779 ( .D0(n4044), .D1(n4045), .D2(n4046), .D3(n4047), .S0(n3756), 
        .S1(n3663), .Y(n4043) );
  MUX4XL U2780 ( .D0(n4034), .D1(n4035), .D2(n4036), .D3(n4037), .S0(n3759), 
        .S1(n3663), .Y(n4023) );
  MUX4XL U2781 ( .D0(n4013), .D1(n4014), .D2(n4015), .D3(n4016), .S0(n3767), 
        .S1(n3664), .Y(n4012) );
  MUX4XL U2782 ( .D0(A[138]), .D1(A[650]), .D2(A[394]), .D3(A[906]), .S0(n3610), .S1(n3700), .Y(n4159) );
  MUX4XL U2783 ( .D0(A[140]), .D1(A[652]), .D2(A[396]), .D3(A[908]), .S0(n3753), .S1(n3694), .Y(n4018) );
  MUX2IXL U2784 ( .D0(n3938), .D1(n3939), .S(n3673), .Y(n3913) );
  MUX2IXL U2785 ( .D0(n3936), .D1(n3937), .S(n3610), .Y(n3935) );
  INVXL U2786 ( .A(n3749), .Y(n3708) );
  MUX2IXL U2787 ( .D0(A[189]), .D1(A[445]), .S(n3693), .Y(n3936) );
  MUX2IXL U2788 ( .D0(A[187]), .D1(A[443]), .S(n3748), .Y(n4077) );
  MUX2IXL U2789 ( .D0(A[185]), .D1(A[441]), .S(n3686), .Y(n4218) );
  MUX2IXL U2790 ( .D0(A[525]), .D1(A[781]), .S(n3689), .Y(n3983) );
  MUX2IXL U2791 ( .D0(A[124]), .D1(A[380]), .S(n3689), .Y(n4027) );
  MUX2IXL U2792 ( .D0(A[132]), .D1(A[388]), .S(n3689), .Y(n4019) );
  MUX2IXL U2793 ( .D0(A[228]), .D1(A[484]), .S(n3689), .Y(n3994) );
  MUX2IXL U2794 ( .D0(A[668]), .D1(A[924]), .S(n3689), .Y(n4016) );
  MUX2X1 U2795 ( .D0(n3769), .D1(n3770), .S(SH[7]), .Y(B[7]) );
  MUX4X1 U2796 ( .D0(n3771), .D1(n3772), .D2(n3773), .D3(n3774), .S0(n3677), 
        .S1(n3682), .Y(n3770) );
  MUX2IX1 U2797 ( .D0(n3775), .D1(n3776), .S(n3672), .Y(n3774) );
  MUX2IX1 U2798 ( .D0(n3777), .D1(n3778), .S(n3659), .Y(n3776) );
  MUX4X1 U2799 ( .D0(A[255]), .D1(A[767]), .D2(A[511]), .D3(A[1023]), .S0(
        n3753), .S1(n3697), .Y(n3778) );
  MUX4X1 U2800 ( .D0(A[247]), .D1(A[759]), .D2(A[503]), .D3(A[1015]), .S0(
        n3760), .S1(n3695), .Y(n3777) );
  MUX4X1 U2801 ( .D0(n3779), .D1(n3780), .D2(n3781), .D3(n3782), .S0(n3658), 
        .S1(n3602), .Y(n3775) );
  NOR2X1 U2802 ( .A(A[999]), .B(n3737), .Y(n3781) );
  MUX2IX1 U2803 ( .D0(A[239]), .D1(A[495]), .S(n3690), .Y(n3780) );
  MUX2IX1 U2804 ( .D0(A[231]), .D1(A[487]), .S(n3690), .Y(n3779) );
  MUX4X1 U2805 ( .D0(n3783), .D1(n3784), .D2(n3785), .D3(n3786), .S0(n3671), 
        .S1(n3665), .Y(n3773) );
  MUX2IX1 U2806 ( .D0(n3787), .D1(n3788), .S(n3753), .Y(n3786) );
  NOR2X1 U2807 ( .A(A[991]), .B(n3739), .Y(n3788) );
  NAND2X1 U2808 ( .A(n3789), .B(n3758), .Y(n3785) );
  MUX2IX1 U2809 ( .D0(A[719]), .D1(A[975]), .S(n3691), .Y(n3789) );
  NAND31X1 U2810 ( .C(A[983]), .A(n3700), .B(n3762), .Y(n3784) );
  NAND31X1 U2811 ( .C(A[967]), .A(n3700), .B(n3762), .Y(n3783) );
  MUX4X1 U2812 ( .D0(n3790), .D1(n3791), .D2(n3792), .D3(n3793), .S0(n3671), 
        .S1(n3666), .Y(n3772) );
  MUX2IX1 U2813 ( .D0(n3794), .D1(n3795), .S(n3653), .Y(n3793) );
  NOR2X1 U2814 ( .A(n3703), .B(A[703]), .Y(n3795) );
  MUX2IX1 U2815 ( .D0(A[191]), .D1(A[447]), .S(n3691), .Y(n3794) );
  MUX4X1 U2816 ( .D0(A[175]), .D1(A[687]), .D2(A[431]), .D3(A[943]), .S0(n3753), .S1(n3696), .Y(n3792) );
  MUX4X1 U2817 ( .D0(A[183]), .D1(A[695]), .D2(A[439]), .D3(A[951]), .S0(n3760), .S1(n3696), .Y(n3791) );
  MUX4X1 U2818 ( .D0(A[167]), .D1(A[679]), .D2(A[423]), .D3(A[935]), .S0(n3753), .S1(n3696), .Y(n3790) );
  MUX2IX1 U2819 ( .D0(n3796), .D1(n3797), .S(n3673), .Y(n3771) );
  MUX4X1 U2820 ( .D0(n3798), .D1(n3799), .D2(n3800), .D3(n3801), .S0(n3606), 
        .S1(n3667), .Y(n3797) );
  MUX2IX1 U2821 ( .D0(A[671]), .D1(A[927]), .S(n3691), .Y(n3801) );
  NOR2X1 U2822 ( .A(A[415]), .B(n3738), .Y(n3800) );
  MUX2IX1 U2823 ( .D0(A[663]), .D1(A[919]), .S(n3691), .Y(n3799) );
  NOR2X1 U2824 ( .A(A[407]), .B(n3739), .Y(n3798) );
  MUX2IX1 U2825 ( .D0(n3802), .D1(n3803), .S(n3662), .Y(n3796) );
  MUX4X1 U2826 ( .D0(A[143]), .D1(A[655]), .D2(A[399]), .D3(A[911]), .S0(n3624), .S1(n3697), .Y(n3803) );
  NAND2X1 U2827 ( .A(n3804), .B(n3634), .Y(n3802) );
  MUX2IX1 U2828 ( .D0(A[135]), .D1(A[391]), .S(n3691), .Y(n3804) );
  MUX2IX1 U2829 ( .D0(n3805), .D1(n3806), .S(n3681), .Y(n3769) );
  MUX4X1 U2830 ( .D0(n3807), .D1(n3808), .D2(n3809), .D3(n3810), .S0(n3677), 
        .S1(n3674), .Y(n3806) );
  NOR2X1 U2831 ( .A(n3701), .B(A[639]), .Y(n3814) );
  NOR2X1 U2832 ( .A(n3702), .B(A[631]), .Y(n3813) );
  MUX2IX1 U2833 ( .D0(A[127]), .D1(A[383]), .S(n3693), .Y(n3812) );
  NOR2X1 U2834 ( .A(A[375]), .B(n3738), .Y(n3811) );
  MUX2IX1 U2835 ( .D0(n3815), .D1(n3816), .S(n3662), .Y(n3809) );
  MUX2IX1 U2836 ( .D0(n3817), .D1(n3818), .S(n3759), .Y(n3816) );
  NOR2X1 U2837 ( .A(n3701), .B(A[607]), .Y(n3818) );
  NOR2X1 U2838 ( .A(A[351]), .B(n3737), .Y(n3817) );
  NAND32X1 U2839 ( .B(A[599]), .C(n3743), .A(n3763), .Y(n3815) );
  MUX4X1 U2840 ( .D0(n3819), .D1(n3820), .D2(n3821), .D3(n3822), .S0(n3604), 
        .S1(n3666), .Y(n3808) );
  NOR2X1 U2841 ( .A(n3701), .B(A[623]), .Y(n3822) );
  NOR2X1 U2842 ( .A(A[367]), .B(n3738), .Y(n3821) );
  NOR2X1 U2843 ( .A(n3702), .B(A[615]), .Y(n3820) );
  NOR2X1 U2844 ( .A(A[359]), .B(n3737), .Y(n3819) );
  MUX2X1 U2845 ( .D0(n3823), .D1(n3824), .S(n3667), .Y(n3807) );
  NOR3XL U2846 ( .A(n3634), .B(A[839]), .C(n3706), .Y(n3823) );
  MUX4X1 U2847 ( .D0(n3825), .D1(n3826), .D2(n3827), .D3(n3828), .S0(n3677), 
        .S1(n3675), .Y(n3805) );
  MUX4X1 U2848 ( .D0(n3829), .D1(n3830), .D2(n3831), .D3(n3832), .S0(n3759), 
        .S1(n3666), .Y(n3828) );
  MUX2IX1 U2849 ( .D0(A[575]), .D1(A[831]), .S(n3691), .Y(n3832) );
  NOR2X1 U2850 ( .A(A[319]), .B(n3733), .Y(n3831) );
  MUX2IX1 U2851 ( .D0(A[567]), .D1(A[823]), .S(n3691), .Y(n3830) );
  NOR2X1 U2852 ( .A(A[311]), .B(n3738), .Y(n3829) );
  MUX4X1 U2853 ( .D0(n3833), .D1(n3834), .D2(n3835), .D3(n3836), .S0(n3758), 
        .S1(n3666), .Y(n3827) );
  MUX2IX1 U2854 ( .D0(A[543]), .D1(A[799]), .S(n3691), .Y(n3836) );
  MUX2IX1 U2855 ( .D0(A[535]), .D1(A[791]), .S(n3691), .Y(n3834) );
  NOR2X1 U2856 ( .A(A[279]), .B(n3737), .Y(n3833) );
  MUX2IX1 U2857 ( .D0(n3837), .D1(n3838), .S(n3662), .Y(n3826) );
  MUX4X1 U2858 ( .D0(A[47]), .D1(A[559]), .D2(A[303]), .D3(A[815]), .S0(n3759), 
        .S1(n3699), .Y(n3838) );
  MUX4X1 U2859 ( .D0(A[39]), .D1(A[551]), .D2(A[295]), .D3(A[807]), .S0(n3767), 
        .S1(n3700), .Y(n3837) );
  NOR2X1 U2860 ( .A(n3670), .B(n3839), .Y(n3825) );
  MUX2IX1 U2861 ( .D0(n3840), .D1(n3841), .S(n3753), .Y(n3839) );
  MUX2IX1 U2862 ( .D0(A[527]), .D1(A[783]), .S(n3692), .Y(n3841) );
  NOR2X1 U2863 ( .A(A[271]), .B(n3736), .Y(n3840) );
  MUX2X1 U2864 ( .D0(n3842), .D1(n3843), .S(SH[7]), .Y(B[6]) );
  MUX4X1 U2865 ( .D0(n3844), .D1(n3845), .D2(n3846), .D3(n3847), .S0(n3677), 
        .S1(n3682), .Y(n3843) );
  MUX2IX1 U2866 ( .D0(n3848), .D1(n3849), .S(n3672), .Y(n3847) );
  MUX2IX1 U2867 ( .D0(n3850), .D1(n3851), .S(n3662), .Y(n3849) );
  MUX4X1 U2868 ( .D0(A[246]), .D1(A[758]), .D2(A[502]), .D3(A[1014]), .S0(
        n3756), .S1(n3699), .Y(n3850) );
  MUX4X1 U2869 ( .D0(n3852), .D1(n3853), .D2(n3854), .D3(n3855), .S0(n3658), 
        .S1(n3766), .Y(n3848) );
  NOR2X1 U2870 ( .A(A[1006]), .B(n3732), .Y(n3855) );
  NOR2X1 U2871 ( .A(A[998]), .B(n3736), .Y(n3854) );
  MUX2IX1 U2872 ( .D0(A[238]), .D1(A[494]), .S(n3692), .Y(n3853) );
  MUX2IX1 U2873 ( .D0(A[230]), .D1(A[486]), .S(n3692), .Y(n3852) );
  MUX4X1 U2874 ( .D0(n3856), .D1(n3857), .D2(n3858), .D3(n3859), .S0(n3671), 
        .S1(n3665), .Y(n3846) );
  MUX2IX1 U2875 ( .D0(n3860), .D1(n3861), .S(n3610), .Y(n3859) );
  NOR2X1 U2876 ( .A(A[990]), .B(n3736), .Y(n3861) );
  NAND2X1 U2877 ( .A(n3862), .B(n3604), .Y(n3858) );
  NAND31X1 U2878 ( .C(A[982]), .A(n3748), .B(n3762), .Y(n3857) );
  NAND31X1 U2879 ( .C(A[966]), .A(n3741), .B(n3762), .Y(n3856) );
  NOR2X1 U2880 ( .A(n3750), .B(A[702]), .Y(n3868) );
  MUX2IX1 U2881 ( .D0(A[190]), .D1(A[446]), .S(n3692), .Y(n3867) );
  MUX4X1 U2882 ( .D0(A[174]), .D1(A[686]), .D2(A[430]), .D3(A[942]), .S0(n3604), .S1(n3698), .Y(n3865) );
  MUX4X1 U2883 ( .D0(A[182]), .D1(A[694]), .D2(A[438]), .D3(A[950]), .S0(n3761), .S1(n3698), .Y(n3864) );
  MUX4X1 U2884 ( .D0(A[166]), .D1(A[678]), .D2(A[422]), .D3(A[934]), .S0(n3624), .S1(n3698), .Y(n3863) );
  MUX2IX1 U2885 ( .D0(n3869), .D1(n3870), .S(n3673), .Y(n3844) );
  MUX4X1 U2886 ( .D0(n3871), .D1(n3872), .D2(n3873), .D3(n3874), .S0(n3756), 
        .S1(n3665), .Y(n3870) );
  MUX2IX1 U2887 ( .D0(A[670]), .D1(A[926]), .S(n3692), .Y(n3874) );
  NOR2X1 U2888 ( .A(A[414]), .B(n3735), .Y(n3873) );
  MUX2IX1 U2889 ( .D0(A[662]), .D1(A[918]), .S(n3692), .Y(n3872) );
  NOR2X1 U2890 ( .A(A[406]), .B(n3736), .Y(n3871) );
  MUX2IX1 U2891 ( .D0(n3875), .D1(n3876), .S(n3662), .Y(n3869) );
  MUX4X1 U2892 ( .D0(A[142]), .D1(A[654]), .D2(A[398]), .D3(A[910]), .S0(n3610), .S1(n3698), .Y(n3876) );
  NAND2X1 U2893 ( .A(n3877), .B(n3765), .Y(n3875) );
  MUX2IX1 U2894 ( .D0(A[134]), .D1(A[390]), .S(n3692), .Y(n3877) );
  MUX2IX1 U2895 ( .D0(n3878), .D1(n3879), .S(n3681), .Y(n3842) );
  MUX4X1 U2896 ( .D0(n3880), .D1(n3881), .D2(n3882), .D3(n3883), .S0(n3677), 
        .S1(n3675), .Y(n3879) );
  MUX4X1 U2897 ( .D0(n3884), .D1(n3885), .D2(n3886), .D3(n3887), .S0(n3658), 
        .S1(n3602), .Y(n3883) );
  NOR2X1 U2898 ( .A(n3702), .B(A[638]), .Y(n3887) );
  NOR2X1 U2899 ( .A(n3702), .B(A[630]), .Y(n3886) );
  MUX2IX1 U2900 ( .D0(A[126]), .D1(A[382]), .S(n3692), .Y(n3885) );
  NOR2X1 U2901 ( .A(A[374]), .B(n3735), .Y(n3884) );
  MUX2IX1 U2902 ( .D0(n3888), .D1(n3889), .S(n3662), .Y(n3882) );
  MUX2IX1 U2903 ( .D0(n3890), .D1(n3891), .S(n3767), .Y(n3889) );
  NOR2X1 U2904 ( .A(n3702), .B(A[606]), .Y(n3891) );
  NOR2X1 U2905 ( .A(A[350]), .B(n3735), .Y(n3890) );
  NAND32X1 U2906 ( .B(A[598]), .C(n3748), .A(n3763), .Y(n3888) );
  MUX4X1 U2907 ( .D0(n3892), .D1(n3740), .D2(n3893), .D3(n3894), .S0(n3659), 
        .S1(n3602), .Y(n3881) );
  NOR2X1 U2908 ( .A(n3703), .B(A[622]), .Y(n3894) );
  NOR2X1 U2909 ( .A(n3703), .B(A[614]), .Y(n3893) );
  NOR2X1 U2910 ( .A(A[358]), .B(n3735), .Y(n3892) );
  MUX2X1 U2911 ( .D0(n3895), .D1(n3824), .S(n3667), .Y(n3880) );
  NOR2X1 U2912 ( .A(n3703), .B(n3764), .Y(n3824) );
  NOR3XL U2913 ( .A(n3764), .B(A[838]), .C(n3727), .Y(n3895) );
  MUX4X1 U2914 ( .D0(n3896), .D1(n3897), .D2(n3898), .D3(n3899), .S0(n3677), 
        .S1(n3675), .Y(n3878) );
  MUX2IX1 U2915 ( .D0(A[574]), .D1(A[830]), .S(n3693), .Y(n3903) );
  NOR2X1 U2916 ( .A(A[318]), .B(n3730), .Y(n3902) );
  MUX2IX1 U2917 ( .D0(A[566]), .D1(A[822]), .S(n3693), .Y(n3901) );
  MUX4X1 U2918 ( .D0(n3904), .D1(n3905), .D2(n3906), .D3(n3907), .S0(n3758), 
        .S1(n3664), .Y(n3898) );
  MUX2IX1 U2919 ( .D0(A[542]), .D1(A[798]), .S(n3693), .Y(n3907) );
  MUX2IX1 U2920 ( .D0(A[534]), .D1(A[790]), .S(n3693), .Y(n3905) );
  NOR2X1 U2921 ( .A(A[278]), .B(n3733), .Y(n3904) );
  MUX2IX1 U2922 ( .D0(n3908), .D1(n3909), .S(n3662), .Y(n3897) );
  MUX4X1 U2923 ( .D0(A[46]), .D1(A[558]), .D2(A[302]), .D3(A[814]), .S0(n3767), 
        .S1(n3694), .Y(n3909) );
  MUX4X1 U2924 ( .D0(A[38]), .D1(A[550]), .D2(A[294]), .D3(A[806]), .S0(n3758), 
        .S1(n3695), .Y(n3908) );
  NOR2X1 U2925 ( .A(n3668), .B(n3910), .Y(n3896) );
  MUX2IX1 U2926 ( .D0(n3911), .D1(n3912), .S(n3756), .Y(n3910) );
  MUX2IX1 U2927 ( .D0(A[526]), .D1(A[782]), .S(n3693), .Y(n3912) );
  NOR2X1 U2928 ( .A(A[270]), .B(n3734), .Y(n3911) );
  MUX2IX1 U2929 ( .D0(n3917), .D1(n3918), .S(n3672), .Y(n3916) );
  MUX2IX1 U2930 ( .D0(n3919), .D1(n3920), .S(n3661), .Y(n3918) );
  MUX4X1 U2931 ( .D0(A[253]), .D1(A[765]), .D2(A[509]), .D3(A[1021]), .S0(
        n3603), .S1(n3694), .Y(n3920) );
  MUX4X1 U2932 ( .D0(A[245]), .D1(A[757]), .D2(A[501]), .D3(A[1013]), .S0(
        n3758), .S1(n3695), .Y(n3919) );
  MUX4X1 U2933 ( .D0(n3921), .D1(n3922), .D2(n3923), .D3(n3924), .S0(n3659), 
        .S1(n3624), .Y(n3917) );
  NOR2X1 U2934 ( .A(A[1005]), .B(n3730), .Y(n3924) );
  NOR2X1 U2935 ( .A(A[997]), .B(n3733), .Y(n3923) );
  MUX2IX1 U2936 ( .D0(A[237]), .D1(A[493]), .S(n3693), .Y(n3922) );
  MUX2IX1 U2937 ( .D0(A[229]), .D1(A[485]), .S(n3694), .Y(n3921) );
  MUX4X1 U2938 ( .D0(n3925), .D1(n3926), .D2(n3927), .D3(n3928), .S0(n3671), 
        .S1(n3664), .Y(n3915) );
  NOR2X1 U2939 ( .A(A[989]), .B(n3732), .Y(n3930) );
  NAND2X1 U2940 ( .A(n3931), .B(n3624), .Y(n3927) );
  NAND31X1 U2941 ( .C(A[965]), .A(n3743), .B(n3753), .Y(n3925) );
  MUX4X1 U2942 ( .D0(n3932), .D1(n3933), .D2(n3934), .D3(n3935), .S0(n3671), 
        .S1(n3664), .Y(n3914) );
  NOR2X1 U2943 ( .A(n3741), .B(A[701]), .Y(n3937) );
  MUX4X1 U2944 ( .D0(A[173]), .D1(A[685]), .D2(A[429]), .D3(A[941]), .S0(n3648), .S1(n3699), .Y(n3934) );
  MUX4X1 U2945 ( .D0(A[165]), .D1(A[677]), .D2(A[421]), .D3(A[933]), .S0(n3766), .S1(n3695), .Y(n3932) );
  MUX4X1 U2946 ( .D0(n3940), .D1(n3941), .D2(n3942), .D3(n3943), .S0(n3606), 
        .S1(n3663), .Y(n3939) );
  MUX2IX1 U2947 ( .D0(A[669]), .D1(A[925]), .S(n3693), .Y(n3943) );
  NOR2X1 U2948 ( .A(A[413]), .B(n3733), .Y(n3942) );
  MUX2IX1 U2949 ( .D0(A[661]), .D1(A[917]), .S(n3690), .Y(n3941) );
  NOR2X1 U2950 ( .A(A[405]), .B(n3732), .Y(n3940) );
  MUX2IX1 U2951 ( .D0(n3944), .D1(n3945), .S(n3662), .Y(n3938) );
  MUX4X1 U2952 ( .D0(A[141]), .D1(A[653]), .D2(A[397]), .D3(A[909]), .S0(n3602), .S1(n3694), .Y(n3945) );
  NAND2X1 U2953 ( .A(n3946), .B(n3764), .Y(n3944) );
  MUX2IX1 U2954 ( .D0(A[133]), .D1(A[389]), .S(n3690), .Y(n3946) );
  MUX4X1 U2955 ( .D0(n3949), .D1(n3950), .D2(n3951), .D3(n3952), .S0(n3677), 
        .S1(n3675), .Y(n3948) );
  MUX4X1 U2956 ( .D0(n3953), .D1(n3954), .D2(n3955), .D3(n3956), .S0(n3659), 
        .S1(n3763), .Y(n3952) );
  NOR2X1 U2957 ( .A(n3740), .B(A[637]), .Y(n3956) );
  NOR2X1 U2958 ( .A(n3703), .B(A[629]), .Y(n3955) );
  MUX2IX1 U2959 ( .D0(A[125]), .D1(A[381]), .S(n3690), .Y(n3954) );
  NOR2X1 U2960 ( .A(A[373]), .B(n3731), .Y(n3953) );
  MUX2IX1 U2961 ( .D0(n3957), .D1(n3958), .S(n3662), .Y(n3951) );
  MUX2IX1 U2962 ( .D0(n3959), .D1(n3960), .S(n3653), .Y(n3958) );
  NOR2X1 U2963 ( .A(n3702), .B(A[605]), .Y(n3960) );
  NOR2X1 U2964 ( .A(A[349]), .B(n3732), .Y(n3959) );
  NAND32X1 U2965 ( .B(A[597]), .C(n3748), .A(n3763), .Y(n3957) );
  MUX4X1 U2966 ( .D0(n3961), .D1(n3962), .D2(n3963), .D3(n3964), .S0(n3606), 
        .S1(n3663), .Y(n3950) );
  NOR2X1 U2967 ( .A(n3702), .B(A[621]), .Y(n3964) );
  NOR2X1 U2968 ( .A(A[365]), .B(n3731), .Y(n3963) );
  NOR2X1 U2969 ( .A(n3742), .B(A[613]), .Y(n3962) );
  NOR2X1 U2970 ( .A(A[357]), .B(n3731), .Y(n3961) );
  MUX2X1 U2971 ( .D0(n3965), .D1(n3966), .S(n3667), .Y(n3949) );
  NOR3XL U2972 ( .A(n3634), .B(n3704), .C(A[589]), .Y(n3966) );
  NOR3XL U2973 ( .A(n3764), .B(A[837]), .C(n3706), .Y(n3965) );
  MUX4X1 U2974 ( .D0(n3967), .D1(n3968), .D2(n3969), .D3(n3970), .S0(n3677), 
        .S1(n3675), .Y(n3947) );
  MUX4X1 U2975 ( .D0(n3971), .D1(n3972), .D2(n3973), .D3(n3974), .S0(n3648), 
        .S1(n3662), .Y(n3970) );
  MUX2IX1 U2976 ( .D0(A[573]), .D1(A[829]), .S(n3690), .Y(n3974) );
  NOR2X1 U2977 ( .A(A[317]), .B(n3731), .Y(n3973) );
  MUX2IX1 U2978 ( .D0(A[565]), .D1(A[821]), .S(n3690), .Y(n3972) );
  NOR2X1 U2979 ( .A(A[309]), .B(n3730), .Y(n3971) );
  MUX4X1 U2980 ( .D0(n3975), .D1(n3976), .D2(n3977), .D3(n3978), .S0(n3759), 
        .S1(n3663), .Y(n3969) );
  MUX2IX1 U2981 ( .D0(A[541]), .D1(A[797]), .S(n3690), .Y(n3978) );
  NOR2X1 U2982 ( .A(A[285]), .B(n3730), .Y(n3977) );
  MUX2IX1 U2983 ( .D0(A[533]), .D1(A[789]), .S(n3690), .Y(n3976) );
  NOR2X1 U2984 ( .A(A[277]), .B(n3729), .Y(n3975) );
  MUX2IX1 U2985 ( .D0(n3979), .D1(n3980), .S(n3661), .Y(n3968) );
  MUX4X1 U2986 ( .D0(A[45]), .D1(A[557]), .D2(A[301]), .D3(A[813]), .S0(n3610), 
        .S1(n3700), .Y(n3980) );
  MUX4X1 U2987 ( .D0(A[37]), .D1(A[549]), .D2(A[293]), .D3(A[805]), .S0(n3604), 
        .S1(n3699), .Y(n3979) );
  NOR2X1 U2988 ( .A(n3668), .B(n3981), .Y(n3967) );
  MUX2IX1 U2989 ( .D0(n3982), .D1(n3983), .S(n3653), .Y(n3981) );
  NOR2X1 U2990 ( .A(A[269]), .B(n3728), .Y(n3982) );
  MUX4X1 U2991 ( .D0(n3986), .D1(n3987), .D2(n3988), .D3(n3989), .S0(n3677), 
        .S1(n3681), .Y(n3985) );
  MUX2IX1 U2992 ( .D0(n3990), .D1(n3991), .S(n3673), .Y(n3989) );
  MUX4X1 U2993 ( .D0(n3994), .D1(n3995), .D2(n3996), .D3(n3997), .S0(n3659), 
        .S1(n3766), .Y(n3990) );
  NOR2X1 U2994 ( .A(A[1004]), .B(n3729), .Y(n3997) );
  NOR2X1 U2995 ( .A(A[996]), .B(n3729), .Y(n3996) );
  MUX2IX1 U2996 ( .D0(A[236]), .D1(A[492]), .S(n3689), .Y(n3995) );
  MUX4X1 U2997 ( .D0(n3998), .D1(n3999), .D2(n4000), .D3(n4001), .S0(n3671), 
        .S1(n3663), .Y(n3988) );
  NOR2X1 U2998 ( .A(A[988]), .B(n3728), .Y(n4003) );
  MUX2IX1 U2999 ( .D0(A[220]), .D1(A[476]), .S(n3689), .Y(n4002) );
  NAND2X1 U3000 ( .A(n4004), .B(n3758), .Y(n4000) );
  MUX2IX1 U3001 ( .D0(A[716]), .D1(A[972]), .S(n3689), .Y(n4004) );
  NAND31X1 U3002 ( .C(A[980]), .A(n3740), .B(n3762), .Y(n3999) );
  NAND31X1 U3003 ( .C(A[964]), .A(n3741), .B(n3767), .Y(n3998) );
  MUX4X1 U3004 ( .D0(n4005), .D1(n4006), .D2(n4007), .D3(n4008), .S0(n3671), 
        .S1(n3663), .Y(n3987) );
  NOR2X1 U3005 ( .A(n3703), .B(A[700]), .Y(n4010) );
  MUX2IX1 U3006 ( .D0(A[188]), .D1(A[444]), .S(n3689), .Y(n4009) );
  MUX4X1 U3007 ( .D0(A[180]), .D1(A[692]), .D2(A[436]), .D3(A[948]), .S0(n3602), .S1(n3694), .Y(n4006) );
  MUX2IX1 U3008 ( .D0(n4011), .D1(n4012), .S(n3673), .Y(n3986) );
  NOR2X1 U3009 ( .A(A[412]), .B(n3729), .Y(n4015) );
  MUX2IX1 U3010 ( .D0(A[660]), .D1(A[916]), .S(n3689), .Y(n4014) );
  NOR2X1 U3011 ( .A(A[404]), .B(n3728), .Y(n4013) );
  MUX2IX1 U3012 ( .D0(n4017), .D1(n4018), .S(n3661), .Y(n4011) );
  NAND2X1 U3013 ( .A(n4019), .B(n3764), .Y(n4017) );
  MUX2IX1 U3014 ( .D0(n4020), .D1(n4021), .S(n3681), .Y(n3984) );
  MUX4X1 U3015 ( .D0(n4022), .D1(n4023), .D2(n4024), .D3(n4025), .S0(n3678), 
        .S1(n3675), .Y(n4021) );
  MUX4X1 U3016 ( .D0(n4026), .D1(n4027), .D2(n4028), .D3(n4029), .S0(n3659), 
        .S1(n3611), .Y(n4025) );
  NOR2X1 U3017 ( .A(n3703), .B(A[636]), .Y(n4029) );
  NOR2X1 U3018 ( .A(n3740), .B(A[628]), .Y(n4028) );
  NOR2X1 U3019 ( .A(A[372]), .B(n3727), .Y(n4026) );
  MUX2IX1 U3020 ( .D0(n4030), .D1(n4031), .S(n3661), .Y(n4024) );
  MUX2IX1 U3021 ( .D0(n4032), .D1(n4033), .S(n3653), .Y(n4031) );
  NOR2X1 U3022 ( .A(n3704), .B(A[604]), .Y(n4033) );
  NOR2X1 U3023 ( .A(A[348]), .B(n3728), .Y(n4032) );
  NAND32X1 U3024 ( .B(A[596]), .C(n3740), .A(n3763), .Y(n4030) );
  NOR2X1 U3025 ( .A(n3740), .B(A[620]), .Y(n4037) );
  NOR2X1 U3026 ( .A(A[364]), .B(n3727), .Y(n4036) );
  NOR2X1 U3027 ( .A(n3698), .B(A[612]), .Y(n4035) );
  NOR2X1 U3028 ( .A(A[356]), .B(n3727), .Y(n4034) );
  MUX2X1 U3029 ( .D0(n4038), .D1(n4039), .S(n3667), .Y(n4022) );
  NOR3XL U3030 ( .A(n3634), .B(n3704), .C(A[588]), .Y(n4039) );
  NOR3XL U3031 ( .A(n3765), .B(A[836]), .C(n3727), .Y(n4038) );
  MUX4X1 U3032 ( .D0(n4040), .D1(n4041), .D2(n4042), .D3(n4043), .S0(n3678), 
        .S1(n3675), .Y(n4020) );
  MUX2IX1 U3033 ( .D0(A[572]), .D1(A[828]), .S(n3740), .Y(n4047) );
  NOR2X1 U3034 ( .A(A[316]), .B(n3727), .Y(n4046) );
  MUX2IX1 U3035 ( .D0(A[564]), .D1(A[820]), .S(n3744), .Y(n4045) );
  NOR2X1 U3036 ( .A(A[308]), .B(n3726), .Y(n4044) );
  MUX4X1 U3037 ( .D0(n4048), .D1(n4049), .D2(n4050), .D3(n4051), .S0(n3607), 
        .S1(n3663), .Y(n4042) );
  MUX2IX1 U3038 ( .D0(A[540]), .D1(A[796]), .S(n3746), .Y(n4051) );
  NOR2X1 U3039 ( .A(A[284]), .B(n3726), .Y(n4050) );
  MUX2IX1 U3040 ( .D0(A[532]), .D1(A[788]), .S(n3742), .Y(n4049) );
  NOR2X1 U3041 ( .A(A[276]), .B(n3726), .Y(n4048) );
  MUX2IX1 U3042 ( .D0(n4052), .D1(n4053), .S(n3661), .Y(n4041) );
  MUX4X1 U3043 ( .D0(A[44]), .D1(A[556]), .D2(A[300]), .D3(A[812]), .S0(n3767), 
        .S1(n3695), .Y(n4053) );
  MUX4X1 U3044 ( .D0(A[36]), .D1(A[548]), .D2(A[292]), .D3(A[804]), .S0(n3604), 
        .S1(n3696), .Y(n4052) );
  NOR2X1 U3045 ( .A(n3669), .B(n4054), .Y(n4040) );
  MUX2IX1 U3046 ( .D0(n4055), .D1(n4056), .S(n3603), .Y(n4054) );
  MUX2IX1 U3047 ( .D0(A[524]), .D1(A[780]), .S(n3690), .Y(n4056) );
  NOR2X1 U3048 ( .A(A[268]), .B(n3725), .Y(n4055) );
  MUX2IX1 U3049 ( .D0(n4062), .D1(n4063), .S(n3661), .Y(n4061) );
  MUX4X1 U3050 ( .D0(A[251]), .D1(A[763]), .D2(A[507]), .D3(A[1019]), .S0(
        n3606), .S1(n3696), .Y(n4063) );
  MUX4X1 U3051 ( .D0(A[243]), .D1(A[755]), .D2(A[499]), .D3(A[1011]), .S0(
        n3607), .S1(n3695), .Y(n4062) );
  NOR2X1 U3052 ( .A(A[1003]), .B(n3725), .Y(n4067) );
  NOR2X1 U3053 ( .A(A[995]), .B(n3725), .Y(n4066) );
  MUX2IX1 U3054 ( .D0(A[235]), .D1(A[491]), .S(n3745), .Y(n4065) );
  MUX2IX1 U3055 ( .D0(A[227]), .D1(A[483]), .S(n3750), .Y(n4064) );
  NOR2X1 U3056 ( .A(A[987]), .B(n3725), .Y(n4072) );
  MUX2IX1 U3057 ( .D0(A[219]), .D1(A[475]), .S(n3741), .Y(n4071) );
  NAND31X1 U3058 ( .C(A[979]), .A(n3745), .B(n3761), .Y(n4069) );
  NAND31X1 U3059 ( .C(A[963]), .A(n3750), .B(n3604), .Y(n4068) );
  MUX4X1 U3060 ( .D0(n4073), .D1(n4074), .D2(n4075), .D3(n4076), .S0(n3672), 
        .S1(n3664), .Y(n4058) );
  MUX2IX1 U3061 ( .D0(n4077), .D1(n4078), .S(n3603), .Y(n4076) );
  NOR2X1 U3062 ( .A(n3703), .B(A[699]), .Y(n4078) );
  MUX4X1 U3063 ( .D0(A[171]), .D1(A[683]), .D2(A[427]), .D3(A[939]), .S0(n3611), .S1(n3696), .Y(n4075) );
  MUX4X1 U3064 ( .D0(A[163]), .D1(A[675]), .D2(A[419]), .D3(A[931]), .S0(n3756), .S1(n3697), .Y(n4073) );
  MUX2IX1 U3065 ( .D0(n4079), .D1(n4080), .S(n3673), .Y(n4057) );
  MUX4X1 U3066 ( .D0(n4081), .D1(n4082), .D2(n4083), .D3(n4084), .S0(n3611), 
        .S1(n3663), .Y(n4080) );
  MUX2IX1 U3067 ( .D0(A[667]), .D1(A[923]), .S(n3688), .Y(n4084) );
  NOR2X1 U3068 ( .A(A[411]), .B(n3724), .Y(n4083) );
  MUX2IX1 U3069 ( .D0(A[659]), .D1(A[915]), .S(n3688), .Y(n4082) );
  NOR2X1 U3070 ( .A(A[403]), .B(n3724), .Y(n4081) );
  MUX2IX1 U3071 ( .D0(n4085), .D1(n4086), .S(n3661), .Y(n4079) );
  MUX4X1 U3072 ( .D0(A[139]), .D1(A[651]), .D2(A[395]), .D3(A[907]), .S0(n3756), .S1(n3697), .Y(n4086) );
  NAND2X1 U3073 ( .A(n4087), .B(n3764), .Y(n4085) );
  MUX2IX1 U3074 ( .D0(A[131]), .D1(A[387]), .S(n3688), .Y(n4087) );
  MUX4X1 U3075 ( .D0(n4090), .D1(n4091), .D2(n4092), .D3(n4093), .S0(n3678), 
        .S1(n3675), .Y(n4089) );
  NOR2X1 U3076 ( .A(n3702), .B(A[635]), .Y(n4097) );
  NOR2X1 U3077 ( .A(n3702), .B(A[627]), .Y(n4096) );
  MUX2IX1 U3078 ( .D0(A[123]), .D1(A[379]), .S(n3688), .Y(n4095) );
  NOR2X1 U3079 ( .A(A[371]), .B(n3724), .Y(n4094) );
  MUX2IX1 U3080 ( .D0(n4098), .D1(n4099), .S(n3660), .Y(n4092) );
  MUX2IX1 U3081 ( .D0(n4100), .D1(n4101), .S(n3604), .Y(n4099) );
  NOR2X1 U3082 ( .A(n3701), .B(A[603]), .Y(n4101) );
  NOR2X1 U3083 ( .A(A[347]), .B(n3724), .Y(n4100) );
  NAND32X1 U3084 ( .B(A[595]), .C(n3740), .A(n3763), .Y(n4098) );
  MUX4X1 U3085 ( .D0(n4102), .D1(n4103), .D2(n4104), .D3(n4105), .S0(n3624), 
        .S1(n3664), .Y(n4091) );
  NOR2X1 U3086 ( .A(n3741), .B(A[619]), .Y(n4105) );
  NOR2X1 U3087 ( .A(A[363]), .B(n3723), .Y(n4104) );
  NOR2X1 U3088 ( .A(n3701), .B(A[611]), .Y(n4103) );
  NOR2X1 U3089 ( .A(A[355]), .B(n3723), .Y(n4102) );
  MUX2X1 U3090 ( .D0(n4106), .D1(n4107), .S(n3660), .Y(n4090) );
  NOR3XL U3091 ( .A(n3765), .B(n3704), .C(A[587]), .Y(n4107) );
  NOR3XL U3092 ( .A(n3765), .B(A[835]), .C(n3739), .Y(n4106) );
  MUX4X1 U3093 ( .D0(n4108), .D1(n4109), .D2(n4110), .D3(n4111), .S0(n3678), 
        .S1(n3674), .Y(n4088) );
  MUX4X1 U3094 ( .D0(n4112), .D1(n4113), .D2(n4114), .D3(n4115), .S0(n3759), 
        .S1(n3664), .Y(n4111) );
  MUX2IX1 U3095 ( .D0(A[571]), .D1(A[827]), .S(n3688), .Y(n4115) );
  NOR2X1 U3096 ( .A(A[315]), .B(n3723), .Y(n4114) );
  MUX2IX1 U3097 ( .D0(A[563]), .D1(A[819]), .S(n3688), .Y(n4113) );
  NOR2X1 U3098 ( .A(A[307]), .B(n3723), .Y(n4112) );
  MUX4X1 U3099 ( .D0(n4116), .D1(n4117), .D2(n4118), .D3(n4119), .S0(n3758), 
        .S1(n3664), .Y(n4110) );
  MUX2IX1 U3100 ( .D0(A[539]), .D1(A[795]), .S(n3688), .Y(n4119) );
  NOR2X1 U3101 ( .A(A[283]), .B(n3722), .Y(n4118) );
  MUX2IX1 U3102 ( .D0(A[531]), .D1(A[787]), .S(n3688), .Y(n4117) );
  NOR2X1 U3103 ( .A(A[275]), .B(n3722), .Y(n4116) );
  MUX2IX1 U3104 ( .D0(n4120), .D1(n4121), .S(n3660), .Y(n4109) );
  MUX4X1 U3105 ( .D0(A[43]), .D1(A[555]), .D2(A[299]), .D3(A[811]), .S0(n3653), 
        .S1(n3698), .Y(n4121) );
  MUX4X1 U3106 ( .D0(A[35]), .D1(A[547]), .D2(A[291]), .D3(A[803]), .S0(n3759), 
        .S1(n3698), .Y(n4120) );
  NOR2X1 U3107 ( .A(n3669), .B(n4122), .Y(n4108) );
  MUX2IX1 U3108 ( .D0(n4123), .D1(n4124), .S(n3606), .Y(n4122) );
  MUX2IX1 U3109 ( .D0(A[523]), .D1(A[779]), .S(n3688), .Y(n4124) );
  NOR2X1 U3110 ( .A(A[267]), .B(n3722), .Y(n4123) );
  MUX2X1 U3111 ( .D0(n4125), .D1(n4126), .S(SH[7]), .Y(B[2]) );
  MUX4X1 U3112 ( .D0(n4127), .D1(n4128), .D2(n4129), .D3(n4130), .S0(n3678), 
        .S1(n3682), .Y(n4126) );
  MUX2IX1 U3113 ( .D0(n4131), .D1(n4132), .S(n3674), .Y(n4130) );
  MUX2IX1 U3114 ( .D0(n4133), .D1(n4134), .S(n3661), .Y(n4132) );
  MUX4X1 U3115 ( .D0(A[250]), .D1(A[762]), .D2(A[506]), .D3(A[1018]), .S0(
        n3603), .S1(n3698), .Y(n4134) );
  MUX4X1 U3116 ( .D0(A[242]), .D1(A[754]), .D2(A[498]), .D3(A[1010]), .S0(
        n3648), .S1(n3698), .Y(n4133) );
  MUX4X1 U3117 ( .D0(n4135), .D1(n4136), .D2(n4137), .D3(n4138), .S0(n3659), 
        .S1(n3755), .Y(n4131) );
  NOR2X1 U3118 ( .A(A[1002]), .B(n3722), .Y(n4138) );
  NOR2X1 U3119 ( .A(A[994]), .B(n3721), .Y(n4137) );
  MUX2IX1 U3120 ( .D0(A[234]), .D1(A[490]), .S(n3688), .Y(n4136) );
  MUX2IX1 U3121 ( .D0(A[226]), .D1(A[482]), .S(n3687), .Y(n4135) );
  MUX4X1 U3122 ( .D0(n4139), .D1(n4140), .D2(n4141), .D3(n4142), .S0(n3672), 
        .S1(n3665), .Y(n4129) );
  MUX2IX1 U3123 ( .D0(n4143), .D1(n4144), .S(n3602), .Y(n4142) );
  NOR2X1 U3124 ( .A(A[986]), .B(n3721), .Y(n4144) );
  MUX2IX1 U3125 ( .D0(A[218]), .D1(A[474]), .S(n3687), .Y(n4143) );
  NAND2X1 U3126 ( .A(n4145), .B(n3763), .Y(n4141) );
  NAND31X1 U3127 ( .C(A[978]), .A(n3743), .B(n3762), .Y(n4140) );
  NAND31X1 U3128 ( .C(A[962]), .A(n3747), .B(n3760), .Y(n4139) );
  MUX4X1 U3129 ( .D0(n4146), .D1(n4147), .D2(n4148), .D3(n4149), .S0(n3672), 
        .S1(n3664), .Y(n4128) );
  MUX2IX1 U3130 ( .D0(n4150), .D1(n4151), .S(n3607), .Y(n4149) );
  NOR2X1 U3131 ( .A(n3750), .B(A[698]), .Y(n4151) );
  MUX2IX1 U3132 ( .D0(A[186]), .D1(A[442]), .S(n3687), .Y(n4150) );
  MUX4X1 U3133 ( .D0(A[170]), .D1(A[682]), .D2(A[426]), .D3(A[938]), .S0(n3603), .S1(n3699), .Y(n4148) );
  MUX4X1 U3134 ( .D0(A[178]), .D1(A[690]), .D2(A[434]), .D3(A[946]), .S0(n3606), .S1(n3699), .Y(n4147) );
  MUX4X1 U3135 ( .D0(A[162]), .D1(A[674]), .D2(A[418]), .D3(A[930]), .S0(n3607), .S1(n3699), .Y(n4146) );
  MUX2IX1 U3136 ( .D0(n4152), .D1(n4153), .S(n3674), .Y(n4127) );
  MUX2IX1 U3137 ( .D0(A[666]), .D1(A[922]), .S(n3687), .Y(n4157) );
  NOR2X1 U3138 ( .A(A[410]), .B(n3721), .Y(n4156) );
  MUX2IX1 U3139 ( .D0(A[658]), .D1(A[914]), .S(n3687), .Y(n4155) );
  NOR2X1 U3140 ( .A(A[402]), .B(n3721), .Y(n4154) );
  MUX2IX1 U3141 ( .D0(n4158), .D1(n4159), .S(n3660), .Y(n4152) );
  NAND2X1 U3142 ( .A(n4160), .B(n3634), .Y(n4158) );
  MUX2IX1 U3143 ( .D0(A[130]), .D1(A[386]), .S(n3687), .Y(n4160) );
  MUX4X1 U3144 ( .D0(n4163), .D1(n4164), .D2(n4165), .D3(n4166), .S0(n3678), 
        .S1(n3674), .Y(n4162) );
  MUX4X1 U3145 ( .D0(n4167), .D1(n4168), .D2(n4169), .D3(n4170), .S0(n3659), 
        .S1(n3602), .Y(n4166) );
  NOR2X1 U3146 ( .A(n3750), .B(A[634]), .Y(n4170) );
  NOR2X1 U3147 ( .A(n3701), .B(A[626]), .Y(n4169) );
  MUX2IX1 U3148 ( .D0(A[122]), .D1(A[378]), .S(n3687), .Y(n4168) );
  NOR2X1 U3149 ( .A(A[370]), .B(n3720), .Y(n4167) );
  MUX2IX1 U3150 ( .D0(n4171), .D1(n4172), .S(n3660), .Y(n4165) );
  MUX2IX1 U3151 ( .D0(n4173), .D1(n4174), .S(n3648), .Y(n4172) );
  NOR2X1 U3152 ( .A(n3743), .B(A[602]), .Y(n4174) );
  NOR2X1 U3153 ( .A(A[346]), .B(n3720), .Y(n4173) );
  NAND32X1 U3154 ( .B(A[594]), .C(n3742), .A(n3763), .Y(n4171) );
  NOR2X1 U3155 ( .A(n3741), .B(A[618]), .Y(n4178) );
  NOR2X1 U3156 ( .A(A[362]), .B(n3720), .Y(n4177) );
  NOR2X1 U3157 ( .A(n3750), .B(A[610]), .Y(n4176) );
  NOR2X1 U3158 ( .A(A[354]), .B(n3720), .Y(n4175) );
  MUX2X1 U3159 ( .D0(n4179), .D1(n4180), .S(n3660), .Y(n4163) );
  NOR3XL U3160 ( .A(n3765), .B(n3704), .C(A[586]), .Y(n4180) );
  NOR3XL U3161 ( .A(n3765), .B(A[834]), .C(n3739), .Y(n4179) );
  MUX4X1 U3162 ( .D0(n4181), .D1(n4182), .D2(n4183), .D3(n4184), .S0(n3678), 
        .S1(n3674), .Y(n4161) );
  MUX4X1 U3163 ( .D0(n4185), .D1(n4186), .D2(n4187), .D3(n4188), .S0(n3603), 
        .S1(n3665), .Y(n4184) );
  MUX2IX1 U3164 ( .D0(A[570]), .D1(A[826]), .S(n3687), .Y(n4188) );
  NOR2X1 U3165 ( .A(A[314]), .B(n3719), .Y(n4187) );
  MUX2IX1 U3166 ( .D0(A[562]), .D1(A[818]), .S(n3687), .Y(n4186) );
  NOR2X1 U3167 ( .A(A[306]), .B(n3719), .Y(n4185) );
  MUX4X1 U3168 ( .D0(n4189), .D1(n4190), .D2(n4191), .D3(n4192), .S0(n3603), 
        .S1(n3665), .Y(n4183) );
  MUX2IX1 U3169 ( .D0(A[538]), .D1(A[794]), .S(n3686), .Y(n4192) );
  NOR2X1 U3170 ( .A(A[282]), .B(n3719), .Y(n4191) );
  MUX2IX1 U3171 ( .D0(A[530]), .D1(A[786]), .S(n3686), .Y(n4190) );
  NOR2X1 U3172 ( .A(A[274]), .B(n3719), .Y(n4189) );
  MUX2IX1 U3173 ( .D0(n4193), .D1(n4194), .S(n3660), .Y(n4182) );
  MUX4X1 U3174 ( .D0(A[42]), .D1(A[554]), .D2(A[298]), .D3(A[810]), .S0(n3607), 
        .S1(n3700), .Y(n4194) );
  MUX4X1 U3175 ( .D0(A[34]), .D1(A[546]), .D2(A[290]), .D3(A[802]), .S0(n3756), 
        .S1(n3700), .Y(n4193) );
  NOR2X1 U3176 ( .A(n3668), .B(n4195), .Y(n4181) );
  MUX2IX1 U3177 ( .D0(n4196), .D1(n4197), .S(n3759), .Y(n4195) );
  MUX2IX1 U3178 ( .D0(A[522]), .D1(A[778]), .S(n3686), .Y(n4197) );
  NOR2X1 U3179 ( .A(A[266]), .B(n3718), .Y(n4196) );
  MUX4X1 U3180 ( .D0(A[249]), .D1(A[761]), .D2(A[505]), .D3(A[1017]), .S0(
        n3603), .S1(n3699), .Y(n4202) );
  NOR2X1 U3181 ( .A(A[1001]), .B(n3718), .Y(n4206) );
  NOR2X1 U3182 ( .A(A[993]), .B(n3718), .Y(n4205) );
  MUX2IX1 U3183 ( .D0(A[233]), .D1(A[489]), .S(n3686), .Y(n4204) );
  MUX2IX1 U3184 ( .D0(A[225]), .D1(A[481]), .S(n3686), .Y(n4203) );
  MUX2IX1 U3185 ( .D0(n4211), .D1(n4212), .S(n3610), .Y(n4210) );
  NOR2X1 U3186 ( .A(A[985]), .B(n3718), .Y(n4212) );
  MUX2IX1 U3187 ( .D0(A[217]), .D1(A[473]), .S(n3686), .Y(n4211) );
  MUX2IX1 U3188 ( .D0(A[713]), .D1(A[969]), .S(n3686), .Y(n4213) );
  NAND31X1 U3189 ( .C(A[977]), .A(n3746), .B(n3762), .Y(n4208) );
  NAND31X1 U3190 ( .C(A[961]), .A(n3700), .B(n3767), .Y(n4207) );
  MUX2IX1 U3191 ( .D0(n4218), .D1(n4219), .S(n3766), .Y(n4217) );
  NOR2X1 U3192 ( .A(n3742), .B(A[697]), .Y(n4219) );
  MUX4X1 U3193 ( .D0(A[169]), .D1(A[681]), .D2(A[425]), .D3(A[937]), .S0(n3753), .S1(n3697), .Y(n4216) );
  MUX4X1 U3194 ( .D0(A[177]), .D1(A[689]), .D2(A[433]), .D3(A[945]), .S0(n3761), .S1(n3697), .Y(n4215) );
  MUX4X1 U3195 ( .D0(n4222), .D1(n4223), .D2(n4224), .D3(n4225), .S0(n3758), 
        .S1(n3666), .Y(n4221) );
  MUX2IX1 U3196 ( .D0(A[665]), .D1(A[921]), .S(n3686), .Y(n4225) );
  NOR2X1 U3197 ( .A(A[409]), .B(n3717), .Y(n4224) );
  MUX2IX1 U3198 ( .D0(A[657]), .D1(A[913]), .S(n3686), .Y(n4223) );
  NOR2X1 U3199 ( .A(A[401]), .B(n3717), .Y(n4222) );
  NAND2X1 U3200 ( .A(n4227), .B(n3765), .Y(n4226) );
  MUX2IX1 U3201 ( .D0(A[129]), .D1(A[385]), .S(n3685), .Y(n4227) );
  MUX2IX1 U3202 ( .D0(n4228), .D1(n4229), .S(n3681), .Y(n4198) );
  MUX4X1 U3203 ( .D0(n4230), .D1(n4231), .D2(n4232), .D3(n4233), .S0(n3678), 
        .S1(n3674), .Y(n4229) );
  MUX4X1 U3204 ( .D0(n4234), .D1(n4235), .D2(n4236), .D3(n4237), .S0(n3658), 
        .S1(n3604), .Y(n4233) );
  NOR2X1 U3205 ( .A(n3701), .B(A[633]), .Y(n4237) );
  NOR2X1 U3206 ( .A(n3701), .B(A[625]), .Y(n4236) );
  MUX2IX1 U3207 ( .D0(A[121]), .D1(A[377]), .S(n3685), .Y(n4235) );
  NOR2X1 U3208 ( .A(A[369]), .B(n3717), .Y(n4234) );
  MUX2IX1 U3209 ( .D0(n4238), .D1(n4239), .S(n3660), .Y(n4232) );
  MUX2IX1 U3210 ( .D0(n4240), .D1(n4241), .S(n3766), .Y(n4239) );
  NOR2X1 U3211 ( .A(n3701), .B(A[601]), .Y(n4241) );
  NOR2X1 U3212 ( .A(A[345]), .B(n3717), .Y(n4240) );
  NAND32X1 U3213 ( .B(A[593]), .C(n3742), .A(n3763), .Y(n4238) );
  MUX4X1 U3214 ( .D0(n4242), .D1(n4243), .D2(n4244), .D3(n4245), .S0(n3758), 
        .S1(n3666), .Y(n4231) );
  NOR2X1 U3215 ( .A(n3701), .B(A[617]), .Y(n4245) );
  NOR2X1 U3216 ( .A(A[361]), .B(n3716), .Y(n4244) );
  NOR2X1 U3217 ( .A(n3702), .B(A[609]), .Y(n4243) );
  NOR2X1 U3218 ( .A(A[353]), .B(n3716), .Y(n4242) );
  MUX2X1 U3219 ( .D0(n4246), .D1(n4247), .S(n3661), .Y(n4230) );
  NOR3XL U3220 ( .A(n3634), .B(n3704), .C(A[585]), .Y(n4247) );
  NOR3XL U3221 ( .A(n3634), .B(A[833]), .C(n3727), .Y(n4246) );
  MUX4X1 U3222 ( .D0(n4248), .D1(n4249), .D2(n4250), .D3(n4251), .S0(n3679), 
        .S1(n3674), .Y(n4228) );
  MUX4X1 U3223 ( .D0(n4252), .D1(n4253), .D2(n4254), .D3(n4255), .S0(n3758), 
        .S1(n3666), .Y(n4251) );
  MUX2IX1 U3224 ( .D0(A[569]), .D1(A[825]), .S(n3685), .Y(n4255) );
  NOR2X1 U3225 ( .A(A[313]), .B(n3716), .Y(n4254) );
  MUX2IX1 U3226 ( .D0(A[561]), .D1(A[817]), .S(n3685), .Y(n4253) );
  NOR2X1 U3227 ( .A(A[305]), .B(n3716), .Y(n4252) );
  MUX4X1 U3228 ( .D0(n4256), .D1(n4257), .D2(n4258), .D3(n4259), .S0(n3759), 
        .S1(n3666), .Y(n4250) );
  MUX2IX1 U3229 ( .D0(A[537]), .D1(A[793]), .S(n3685), .Y(n4259) );
  NOR2X1 U3230 ( .A(A[281]), .B(n3715), .Y(n4258) );
  MUX2IX1 U3231 ( .D0(A[529]), .D1(A[785]), .S(n3685), .Y(n4257) );
  NOR2X1 U3232 ( .A(A[273]), .B(n3715), .Y(n4256) );
  MUX2IX1 U3233 ( .D0(n4260), .D1(n4261), .S(n3659), .Y(n4249) );
  MUX4X1 U3234 ( .D0(A[41]), .D1(A[553]), .D2(A[297]), .D3(A[809]), .S0(n3760), 
        .S1(n3697), .Y(n4261) );
  MUX4X1 U3235 ( .D0(A[33]), .D1(A[545]), .D2(A[289]), .D3(A[801]), .S0(n3611), 
        .S1(n3697), .Y(n4260) );
  NOR2X1 U3236 ( .A(n3669), .B(n4262), .Y(n4248) );
  MUX2IX1 U3237 ( .D0(A[521]), .D1(A[777]), .S(n3685), .Y(n4264) );
  NOR2X1 U3238 ( .A(A[265]), .B(n3715), .Y(n4263) );
  MUX4X1 U3239 ( .D0(A[248]), .D1(A[760]), .D2(A[504]), .D3(A[1016]), .S0(
        n3756), .S1(n3696), .Y(n4267) );
  MUX4X1 U3240 ( .D0(A[240]), .D1(A[752]), .D2(A[496]), .D3(A[1008]), .S0(
        n3611), .S1(n3697), .Y(n4266) );
  NOR2X1 U3241 ( .A(A[1000]), .B(n3715), .Y(n4271) );
  NOR2X1 U3242 ( .A(A[992]), .B(n3714), .Y(n4270) );
  MUX2IX1 U3243 ( .D0(A[232]), .D1(A[488]), .S(n3685), .Y(n4269) );
  MUX2IX1 U3244 ( .D0(A[224]), .D1(A[480]), .S(n3685), .Y(n4268) );
  MUX2IX1 U3245 ( .D0(n4276), .D1(n4277), .S(n3754), .Y(n4275) );
  NOR2X1 U3246 ( .A(A[984]), .B(n3714), .Y(n4277) );
  MUX2IX1 U3247 ( .D0(A[216]), .D1(A[472]), .S(n3685), .Y(n4276) );
  NAND2X1 U3248 ( .A(n4278), .B(n3767), .Y(n4274) );
  MUX2IX1 U3249 ( .D0(A[712]), .D1(A[968]), .S(n3684), .Y(n4278) );
  NAND31X1 U3250 ( .C(A[976]), .A(n3750), .B(n3762), .Y(n4273) );
  NAND31X1 U3251 ( .C(A[960]), .A(n3700), .B(n3762), .Y(n4272) );
  MUX2IX1 U3252 ( .D0(n4283), .D1(n4284), .S(n3611), .Y(n4282) );
  NOR2X1 U3253 ( .A(n3703), .B(A[696]), .Y(n4284) );
  MUX2IX1 U3254 ( .D0(A[184]), .D1(A[440]), .S(n3684), .Y(n4283) );
  MUX4X1 U3255 ( .D0(A[168]), .D1(A[680]), .D2(A[424]), .D3(A[936]), .S0(n3648), .S1(n3695), .Y(n4281) );
  MUX4X1 U3256 ( .D0(A[176]), .D1(A[688]), .D2(A[432]), .D3(A[944]), .S0(n3606), .S1(n3695), .Y(n4280) );
  MUX4X1 U3257 ( .D0(A[160]), .D1(A[672]), .D2(A[416]), .D3(A[928]), .S0(n3611), .S1(n3696), .Y(n4279) );
  MUX4X1 U3258 ( .D0(n4287), .D1(n4288), .D2(n4289), .D3(n4290), .S0(n3767), 
        .S1(n3667), .Y(n4286) );
  MUX2IX1 U3259 ( .D0(A[664]), .D1(A[920]), .S(n3684), .Y(n4290) );
  NOR2X1 U3260 ( .A(A[408]), .B(n3714), .Y(n4289) );
  MUX2IX1 U3261 ( .D0(A[656]), .D1(A[912]), .S(n3684), .Y(n4288) );
  NOR2X1 U3262 ( .A(A[400]), .B(n3714), .Y(n4287) );
  MUX2IX1 U3263 ( .D0(n4291), .D1(n4292), .S(n3660), .Y(n4285) );
  MUX4X1 U3264 ( .D0(A[136]), .D1(A[648]), .D2(A[392]), .D3(A[904]), .S0(n3604), .S1(n3695), .Y(n4292) );
  MUX2IX1 U3265 ( .D0(n4293), .D1(n4294), .S(n3681), .Y(n4265) );
  MUX4X1 U3266 ( .D0(n4295), .D1(n4296), .D2(n4297), .D3(n4298), .S0(n3679), 
        .S1(n3674), .Y(n4294) );
  NOR2X1 U3267 ( .A(n3697), .B(A[632]), .Y(n4302) );
  NOR2X1 U3268 ( .A(n3703), .B(A[624]), .Y(n4301) );
  MUX2IX1 U3269 ( .D0(A[120]), .D1(A[376]), .S(n3684), .Y(n4300) );
  NOR2X1 U3270 ( .A(A[368]), .B(n3713), .Y(n4299) );
  MUX2IX1 U3271 ( .D0(n4303), .D1(n4304), .S(n3659), .Y(n4297) );
  NOR2X1 U3272 ( .A(n3742), .B(A[600]), .Y(n4306) );
  NOR2X1 U3273 ( .A(A[344]), .B(n3713), .Y(n4305) );
  NAND32X1 U3274 ( .B(A[592]), .C(n3744), .A(n3763), .Y(n4303) );
  MUX4X1 U3275 ( .D0(n4307), .D1(n4308), .D2(n4309), .D3(n4310), .S0(n3603), 
        .S1(n3667), .Y(n4296) );
  NOR2X1 U3276 ( .A(n3740), .B(A[616]), .Y(n4310) );
  NOR2X1 U3277 ( .A(A[360]), .B(n3713), .Y(n4309) );
  NOR2X1 U3278 ( .A(n3704), .B(A[608]), .Y(n4308) );
  NOR2X1 U3279 ( .A(A[352]), .B(n3713), .Y(n4307) );
  MUX2X1 U3280 ( .D0(n4311), .D1(n4312), .S(SH[3]), .Y(n4295) );
  NOR3XL U3281 ( .A(n3765), .B(n3704), .C(A[584]), .Y(n4312) );
  NOR3XL U3282 ( .A(n3765), .B(A[832]), .C(n3727), .Y(n4311) );
  MUX4X1 U3283 ( .D0(n4313), .D1(n4314), .D2(n4315), .D3(n4316), .S0(n3679), 
        .S1(n3674), .Y(n4293) );
  MUX4X1 U3284 ( .D0(n4317), .D1(n4318), .D2(n4319), .D3(n4320), .S0(n3767), 
        .S1(n3667), .Y(n4316) );
  MUX2IX1 U3285 ( .D0(A[568]), .D1(A[824]), .S(n3684), .Y(n4320) );
  NOR2X1 U3286 ( .A(A[312]), .B(n3712), .Y(n4319) );
  MUX2IX1 U3287 ( .D0(A[560]), .D1(A[816]), .S(n3684), .Y(n4318) );
  NOR2X1 U3288 ( .A(A[304]), .B(n3712), .Y(n4317) );
  MUX4X1 U3289 ( .D0(n4321), .D1(n4322), .D2(n4323), .D3(n4324), .S0(n3602), 
        .S1(n3667), .Y(n4315) );
  MUX2IX1 U3290 ( .D0(A[536]), .D1(A[792]), .S(n3684), .Y(n4324) );
  NOR2X1 U3291 ( .A(A[280]), .B(n3712), .Y(n4323) );
  MUX2IX1 U3292 ( .D0(A[528]), .D1(A[784]), .S(n3684), .Y(n4322) );
  NOR2X1 U3293 ( .A(A[272]), .B(n3712), .Y(n4321) );
  MUX2IX1 U3294 ( .D0(n4325), .D1(n4326), .S(n3661), .Y(n4314) );
  MUX4X1 U3295 ( .D0(A[40]), .D1(A[552]), .D2(A[296]), .D3(A[808]), .S0(n3761), 
        .S1(n3695), .Y(n4326) );
  MUX4X1 U3296 ( .D0(A[32]), .D1(A[544]), .D2(A[288]), .D3(A[800]), .S0(n3760), 
        .S1(n3694), .Y(n4325) );
  NOR2X1 U3297 ( .A(n3669), .B(n4327), .Y(n4313) );
  MUX2IX1 U3298 ( .D0(n4328), .D1(n4329), .S(n3759), .Y(n4327) );
  MUX2IX1 U3299 ( .D0(A[520]), .D1(A[776]), .S(n3744), .Y(n4329) );
  NOR2X1 U3300 ( .A(A[264]), .B(n3726), .Y(n4328) );
endmodule


module regbank_a0_DW01_inc_0 ( A, SUM );
  input [15:0] A;
  output [15:0] SUM;

  wire   [14:2] carry;

  HAD1X1 U1_1_13 ( .A(A[13]), .B(carry[13]), .CO(carry[14]), .SO(SUM[13]) );
  HAD1X1 U1_1_12 ( .A(A[12]), .B(carry[12]), .CO(carry[13]), .SO(SUM[12]) );
  HAD1X1 U1_1_11 ( .A(A[11]), .B(carry[11]), .CO(carry[12]), .SO(SUM[11]) );
  HAD1X1 U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .SO(SUM[10]) );
  HAD1X1 U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .SO(SUM[9]) );
  HAD1X1 U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .SO(SUM[8]) );
  HAD1X1 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .SO(SUM[7]) );
  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  XOR2X1 U1_1_14 ( .A(A[14]), .B(carry[14]), .Y(SUM[14]) );
  INVX1 U1 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module regbank_a0_DW01_add_0 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;

  wire   [7:1] carry;

  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  XOR3X1 U1_7 ( .A(A[7]), .B(B[7]), .C(carry[7]), .Y(SUM[7]) );
  AND2X1 U1 ( .A(A[0]), .B(B[0]), .Y(carry[1]) );
  XOR2X1 U2 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_regbank_a0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_49 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net10776;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_49 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10776), .TE(1'b0) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net10776), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net10776), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net10776), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net10776), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net10776), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net10776), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net10776), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net10776), .XR(arstz), .Q(rdat[4]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_49 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_50 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net10794;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_50 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10794), .TE(1'b0) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net10794), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net10794), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net10794), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net10794), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net10794), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net10794), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net10794), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net10794), .XR(arstz), .Q(rdat[4]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_50 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_51 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net10812;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_51 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10812), .TE(1'b0) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net10812), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net10812), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net10812), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net10812), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net10812), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net10812), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net10812), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net10812), .XR(arstz), .Q(rdat[5]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_51 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_52 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net10830;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_52 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10830), .TE(1'b0) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net10830), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net10830), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net10830), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net10830), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net10830), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net10830), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net10830), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net10830), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_52 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_53 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net10848;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_53 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10848), .TE(1'b0) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net10848), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net10848), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net10848), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net10848), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net10848), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net10848), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net10848), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net10848), .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_53 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_8_0000001f ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net10866;

  SNPS_CLOCK_GATE_HIGH_glreg_8_0000001f clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10866), .TE(1'b0) );
  DFFSQX1 mem_reg_3_ ( .D(wdat[3]), .C(net10866), .XS(arstz), .Q(rdat[3]) );
  DFFSQX1 mem_reg_2_ ( .D(wdat[2]), .C(net10866), .XS(arstz), .Q(rdat[2]) );
  DFFSQX1 mem_reg_1_ ( .D(wdat[1]), .C(net10866), .XS(arstz), .Q(rdat[1]) );
  DFFSQX1 mem_reg_0_ ( .D(wdat[0]), .C(net10866), .XS(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net10866), .XR(arstz), .Q(rdat[7]) );
  DFFSQX1 mem_reg_4_ ( .D(wdat[4]), .C(net10866), .XS(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net10866), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net10866), .XR(arstz), .Q(rdat[5]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_8_0000001f ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_8_00000004 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net10884;

  SNPS_CLOCK_GATE_HIGH_glreg_8_00000004 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10884), .TE(1'b0) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net10884), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net10884), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net10884), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net10884), .XR(arstz), .Q(rdat[6]) );
  DFFSQX1 mem_reg_2_ ( .D(wdat[2]), .C(net10884), .XS(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net10884), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net10884), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net10884), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_8_00000004 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_4_00000004 ( clk, arstz, we, wdat, rdat );
  input [3:0] wdat;
  output [3:0] rdat;
  input clk, arstz, we;
  wire   net10902;

  SNPS_CLOCK_GATE_HIGH_glreg_4_00000004 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10902), .TE(1'b0) );
  DFFSQX1 mem_reg_2_ ( .D(wdat[2]), .C(net10902), .XS(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net10902), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net10902), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net10902), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_4_00000004 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_54 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net10920;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_54 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10920), .TE(1'b0) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net10920), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net10920), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net10920), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net10920), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net10920), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net10920), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net10920), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net10920), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_54 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_55 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net10938;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_55 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10938), .TE(1'b0) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net10938), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net10938), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net10938), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net10938), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net10938), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net10938), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net10938), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net10938), .XR(arstz), .Q(rdat[2]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_55 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glsta_a0_2 ( clk, arstz, rst0, set2, clr1, rdat, irq );
  input [7:0] set2;
  input [7:0] clr1;
  output [7:0] rdat;
  output [7:0] irq;
  input clk, arstz, rst0;
  wire   upd_r, n17, n18, n19, n20, n21, n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16;
  wire   [7:0] wd_r;

  glreg_WIDTH8_2 u0 ( .clk(clk), .arstz(arstz), .we(upd_r), .wdat(wd_r), 
        .rdat(rdat) );
  NOR4XL U2 ( .A(clr1[7]), .B(clr1[6]), .C(clr1[5]), .D(clr1[4]), .Y(n18) );
  INVX1 U3 ( .A(set2[2]), .Y(n1) );
  INVX1 U4 ( .A(set2[4]), .Y(n2) );
  INVX1 U5 ( .A(set2[5]), .Y(n3) );
  INVX1 U6 ( .A(set2[7]), .Y(n12) );
  INVX1 U7 ( .A(set2[0]), .Y(n13) );
  INVX1 U8 ( .A(set2[1]), .Y(n14) );
  INVX1 U9 ( .A(set2[3]), .Y(n15) );
  NAND3X1 U10 ( .A(n16), .B(n12), .C(n3), .Y(n21) );
  NAND4X1 U11 ( .A(n17), .B(n18), .C(n19), .D(n20), .Y(upd_r) );
  NOR4XL U12 ( .A(set2[2]), .B(set2[1]), .C(set2[0]), .D(rst0), .Y(n19) );
  NOR3XL U13 ( .A(n21), .B(set2[4]), .C(set2[3]), .Y(n20) );
  NOR4XL U14 ( .A(clr1[3]), .B(clr1[2]), .C(clr1[1]), .D(clr1[0]), .Y(n17) );
  AOI211X1 U15 ( .C(n13), .D(n11), .A(rst0), .B(clr1[0]), .Y(wd_r[0]) );
  INVX1 U16 ( .A(rdat[0]), .Y(n11) );
  AOI211X1 U17 ( .C(n14), .D(n10), .A(rst0), .B(clr1[1]), .Y(wd_r[1]) );
  INVX1 U18 ( .A(rdat[1]), .Y(n10) );
  AOI211X1 U19 ( .C(n1), .D(n9), .A(rst0), .B(clr1[2]), .Y(wd_r[2]) );
  INVX1 U20 ( .A(rdat[2]), .Y(n9) );
  AOI211X1 U21 ( .C(n15), .D(n8), .A(rst0), .B(clr1[3]), .Y(wd_r[3]) );
  INVX1 U22 ( .A(rdat[3]), .Y(n8) );
  AOI211X1 U23 ( .C(n2), .D(n7), .A(rst0), .B(clr1[4]), .Y(wd_r[4]) );
  INVX1 U24 ( .A(rdat[4]), .Y(n7) );
  AOI211X1 U25 ( .C(n3), .D(n6), .A(rst0), .B(clr1[5]), .Y(wd_r[5]) );
  INVX1 U26 ( .A(rdat[5]), .Y(n6) );
  AOI211X1 U27 ( .C(n16), .D(n5), .A(rst0), .B(clr1[6]), .Y(wd_r[6]) );
  INVX1 U28 ( .A(rdat[6]), .Y(n5) );
  AOI211X1 U29 ( .C(n12), .D(n4), .A(rst0), .B(clr1[7]), .Y(wd_r[7]) );
  INVX1 U30 ( .A(rdat[7]), .Y(n4) );
  NOR2X1 U31 ( .A(rdat[3]), .B(n15), .Y(irq[3]) );
  NOR2X1 U32 ( .A(rdat[2]), .B(n1), .Y(irq[2]) );
  NOR2X1 U33 ( .A(rdat[5]), .B(n3), .Y(irq[5]) );
  NOR2X1 U34 ( .A(rdat[4]), .B(n2), .Y(irq[4]) );
  NOR2X1 U35 ( .A(rdat[0]), .B(n13), .Y(irq[0]) );
  NOR2X1 U36 ( .A(rdat[1]), .B(n14), .Y(irq[1]) );
  NOR2X1 U37 ( .A(rdat[7]), .B(n12), .Y(irq[7]) );
  NOR2X1 U38 ( .A(rdat[6]), .B(n16), .Y(irq[6]) );
  INVX1 U39 ( .A(set2[6]), .Y(n16) );
endmodule


module glreg_WIDTH8_2 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net10956;

  SNPS_CLOCK_GATE_HIGH_glreg_WIDTH8_2 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net10956), .TE(1'b0) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net10956), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net10956), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net10956), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net10956), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net10956), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net10956), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net10956), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net10956), .XR(arstz), .Q(rdat[4]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_WIDTH8_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module dbnc_WIDTH2_TIMEOUT2_8 ( o_dbc, o_chg, i_org, clk, rstz );
  input i_org, clk, rstz;
  output o_dbc, o_chg;
  wire   d_org_0_, n1, n7, n8, n9, n10, n11;
  wire   [1:0] db_cnt;

  DFFRQX1 db_cnt_reg_1_ ( .D(n8), .C(clk), .XR(rstz), .Q(db_cnt[1]) );
  DFFRQX1 db_cnt_reg_0_ ( .D(n7), .C(clk), .XR(rstz), .Q(db_cnt[0]) );
  DFFRQX1 d_org_reg_0_ ( .D(i_org), .C(clk), .XR(rstz), .Q(d_org_0_) );
  DFFRQX1 d_org_reg_1_ ( .D(n9), .C(clk), .XR(rstz), .Q(o_dbc) );
  NOR32XL U3 ( .B(n11), .C(db_cnt[1]), .A(db_cnt[0]), .Y(o_chg) );
  XNOR2XL U4 ( .A(n1), .B(d_org_0_), .Y(n11) );
  INVX1 U5 ( .A(o_dbc), .Y(n1) );
  ENOX1 U6 ( .A(o_chg), .B(n1), .C(d_org_0_), .D(o_chg), .Y(n9) );
  NAND21X1 U7 ( .B(db_cnt[1]), .A(n11), .Y(n10) );
  NOR21XL U8 ( .B(db_cnt[0]), .A(n10), .Y(n8) );
  NOR2X1 U9 ( .A(db_cnt[0]), .B(n10), .Y(n7) );
endmodule


module dbnc_WIDTH2_TIMEOUT2_9 ( o_dbc, o_chg, i_org, clk, rstz );
  input i_org, clk, rstz;
  output o_dbc, o_chg;
  wire   d_org_0_, n1, n7, n8, n9, n10, n11;
  wire   [1:0] db_cnt;

  DFFRQX1 db_cnt_reg_1_ ( .D(n8), .C(clk), .XR(rstz), .Q(db_cnt[1]) );
  DFFRQX1 db_cnt_reg_0_ ( .D(n7), .C(clk), .XR(rstz), .Q(db_cnt[0]) );
  DFFRQX1 d_org_reg_0_ ( .D(i_org), .C(clk), .XR(rstz), .Q(d_org_0_) );
  DFFRQX1 d_org_reg_1_ ( .D(n9), .C(clk), .XR(rstz), .Q(o_dbc) );
  NOR32XL U3 ( .B(n11), .C(db_cnt[1]), .A(db_cnt[0]), .Y(o_chg) );
  XNOR2XL U4 ( .A(n1), .B(d_org_0_), .Y(n11) );
  INVX1 U5 ( .A(o_dbc), .Y(n1) );
  ENOX1 U6 ( .A(o_chg), .B(n1), .C(d_org_0_), .D(o_chg), .Y(n9) );
  NAND21X1 U7 ( .B(db_cnt[1]), .A(n11), .Y(n10) );
  NOR21XL U8 ( .B(db_cnt[0]), .A(n10), .Y(n8) );
  NOR2X1 U9 ( .A(db_cnt[0]), .B(n10), .Y(n7) );
endmodule


module dbnc_WIDTH2_TIMEOUT2_10 ( o_dbc, o_chg, i_org, clk, rstz );
  input i_org, clk, rstz;
  output o_dbc, o_chg;
  wire   d_org_0_, n1, n7, n8, n9, n10, n11;
  wire   [1:0] db_cnt;

  DFFRQX1 db_cnt_reg_1_ ( .D(n8), .C(clk), .XR(rstz), .Q(db_cnt[1]) );
  DFFRQX1 db_cnt_reg_0_ ( .D(n7), .C(clk), .XR(rstz), .Q(db_cnt[0]) );
  DFFRQX1 d_org_reg_0_ ( .D(i_org), .C(clk), .XR(rstz), .Q(d_org_0_) );
  DFFRQX1 d_org_reg_1_ ( .D(n9), .C(clk), .XR(rstz), .Q(o_dbc) );
  NOR32XL U3 ( .B(n11), .C(db_cnt[1]), .A(db_cnt[0]), .Y(o_chg) );
  XNOR2XL U4 ( .A(n1), .B(d_org_0_), .Y(n11) );
  INVX1 U5 ( .A(o_dbc), .Y(n1) );
  ENOX1 U6 ( .A(o_chg), .B(n1), .C(d_org_0_), .D(o_chg), .Y(n9) );
  NAND21X1 U7 ( .B(db_cnt[1]), .A(n11), .Y(n10) );
  NOR21XL U8 ( .B(db_cnt[0]), .A(n10), .Y(n8) );
  NOR2X1 U9 ( .A(db_cnt[0]), .B(n10), .Y(n7) );
endmodule


module dbnc_WIDTH2_TIMEOUT2_11 ( o_dbc, o_chg, i_org, clk, rstz );
  input i_org, clk, rstz;
  output o_dbc, o_chg;
  wire   d_org_0_, n1, n7, n8, n9, n10, n11;
  wire   [1:0] db_cnt;

  DFFRQX1 db_cnt_reg_1_ ( .D(n8), .C(clk), .XR(rstz), .Q(db_cnt[1]) );
  DFFRQX1 db_cnt_reg_0_ ( .D(n7), .C(clk), .XR(rstz), .Q(db_cnt[0]) );
  DFFRQX1 d_org_reg_0_ ( .D(i_org), .C(clk), .XR(rstz), .Q(d_org_0_) );
  DFFRQX1 d_org_reg_1_ ( .D(n9), .C(clk), .XR(rstz), .Q(o_dbc) );
  XNOR2XL U3 ( .A(n1), .B(d_org_0_), .Y(n11) );
  ENOX1 U4 ( .A(o_chg), .B(n1), .C(d_org_0_), .D(o_chg), .Y(n9) );
  NOR32XL U5 ( .B(n11), .C(db_cnt[1]), .A(db_cnt[0]), .Y(o_chg) );
  INVX1 U6 ( .A(o_dbc), .Y(n1) );
  NAND21X1 U7 ( .B(db_cnt[1]), .A(n11), .Y(n10) );
  NOR21XL U8 ( .B(db_cnt[0]), .A(n10), .Y(n8) );
  NOR2X1 U9 ( .A(db_cnt[0]), .B(n10), .Y(n7) );
endmodule


module dbnc_WIDTH2_TIMEOUT2_12 ( o_dbc, o_chg, i_org, clk, rstz );
  input i_org, clk, rstz;
  output o_dbc, o_chg;
  wire   d_org_0_, n1, n7, n8, n9, n10, n11;
  wire   [1:0] db_cnt;

  DFFRQX1 db_cnt_reg_1_ ( .D(n8), .C(clk), .XR(rstz), .Q(db_cnt[1]) );
  DFFRQX1 db_cnt_reg_0_ ( .D(n7), .C(clk), .XR(rstz), .Q(db_cnt[0]) );
  DFFRQX1 d_org_reg_0_ ( .D(i_org), .C(clk), .XR(rstz), .Q(d_org_0_) );
  DFFRQX1 d_org_reg_1_ ( .D(n9), .C(clk), .XR(rstz), .Q(o_dbc) );
  XNOR2XL U3 ( .A(n1), .B(d_org_0_), .Y(n11) );
  ENOX1 U4 ( .A(o_chg), .B(n1), .C(d_org_0_), .D(o_chg), .Y(n9) );
  NOR32XL U5 ( .B(n11), .C(db_cnt[1]), .A(db_cnt[0]), .Y(o_chg) );
  INVX1 U6 ( .A(o_dbc), .Y(n1) );
  NAND21X1 U7 ( .B(db_cnt[1]), .A(n11), .Y(n10) );
  NOR21XL U8 ( .B(db_cnt[0]), .A(n10), .Y(n8) );
  NOR2X1 U9 ( .A(db_cnt[0]), .B(n10), .Y(n7) );
endmodule


module dbnc_WIDTH2_TIMEOUT2_13 ( o_dbc, o_chg, i_org, clk, rstz );
  input i_org, clk, rstz;
  output o_dbc, o_chg;
  wire   d_org_0_, n2, n3, n4, n5, n6, n1;
  wire   [1:0] db_cnt;

  DFFRQX1 db_cnt_reg_1_ ( .D(n5), .C(clk), .XR(rstz), .Q(db_cnt[1]) );
  DFFRQX1 db_cnt_reg_0_ ( .D(n6), .C(clk), .XR(rstz), .Q(db_cnt[0]) );
  DFFRQX1 d_org_reg_0_ ( .D(i_org), .C(clk), .XR(rstz), .Q(d_org_0_) );
  DFFRQX1 d_org_reg_1_ ( .D(n4), .C(clk), .XR(rstz), .Q(o_dbc) );
  XNOR2XL U3 ( .A(n1), .B(d_org_0_), .Y(n2) );
  ENOX1 U4 ( .A(o_chg), .B(n1), .C(d_org_0_), .D(o_chg), .Y(n4) );
  NOR32XL U5 ( .B(n2), .C(db_cnt[1]), .A(db_cnt[0]), .Y(o_chg) );
  INVX1 U6 ( .A(o_dbc), .Y(n1) );
  NAND21X1 U7 ( .B(db_cnt[1]), .A(n2), .Y(n3) );
  NOR21XL U8 ( .B(db_cnt[0]), .A(n3), .Y(n5) );
  NOR2X1 U9 ( .A(db_cnt[0]), .B(n3), .Y(n6) );
endmodule


module dbnc_WIDTH3_TIMEOUT5_0 ( o_dbc, o_chg, i_org, clk, rstz );
  input i_org, clk, rstz;
  output o_dbc, o_chg;
  wire   d_org_0_, N13, N14, N15, N16, net10974, n5, n6, n7, n1, n2, n3, n4;
  wire   [2:0] db_cnt;

  SNPS_CLOCK_GATE_HIGH_dbnc_WIDTH3_TIMEOUT5_0 clk_gate_db_cnt_reg ( .CLK(clk), 
        .EN(N13), .ENCLK(net10974), .TE(1'b0) );
  DFFRQX1 db_cnt_reg_2_ ( .D(N16), .C(net10974), .XR(rstz), .Q(db_cnt[2]) );
  DFFRQX1 db_cnt_reg_1_ ( .D(N15), .C(net10974), .XR(rstz), .Q(db_cnt[1]) );
  DFFRQX1 d_org_reg_0_ ( .D(i_org), .C(clk), .XR(rstz), .Q(d_org_0_) );
  DFFRQX1 db_cnt_reg_0_ ( .D(N14), .C(net10974), .XR(rstz), .Q(db_cnt[0]) );
  DFFRQX1 d_org_reg_1_ ( .D(n7), .C(net10974), .XR(rstz), .Q(o_dbc) );
  OAI22X1 U3 ( .A(n4), .B(n1), .C(n6), .D(n3), .Y(N16) );
  INVX1 U4 ( .A(N14), .Y(n1) );
  NAND4X1 U5 ( .A(n5), .B(n2), .C(n3), .D(n4), .Y(N13) );
  XNOR2XL U6 ( .A(o_dbc), .B(d_org_0_), .Y(n5) );
  NOR4XL U7 ( .A(n4), .B(n2), .C(n5), .D(db_cnt[1]), .Y(o_chg) );
  INVX1 U8 ( .A(db_cnt[0]), .Y(n2) );
  AO22AXL U9 ( .A(d_org_0_), .B(o_chg), .C(o_dbc), .D(o_chg), .Y(n7) );
  INVX1 U10 ( .A(db_cnt[2]), .Y(n4) );
  NAND31X1 U11 ( .C(n5), .A(n4), .B(db_cnt[0]), .Y(n6) );
  NOR2X1 U12 ( .A(n5), .B(db_cnt[0]), .Y(N14) );
  OAI22X1 U13 ( .A(n3), .B(n1), .C(db_cnt[1]), .D(n6), .Y(N15) );
  INVX1 U14 ( .A(db_cnt[1]), .Y(n3) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dbnc_WIDTH3_TIMEOUT5_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module dbnc_WIDTH3_TIMEOUT5_1 ( o_dbc, o_chg, i_org, clk, rstz );
  input i_org, clk, rstz;
  output o_dbc, o_chg;
  wire   d_org_0_, N13, N14, N15, N16, net10992, n5, n6, n7, n1, n2, n3, n4;
  wire   [2:0] db_cnt;

  SNPS_CLOCK_GATE_HIGH_dbnc_WIDTH3_TIMEOUT5_1 clk_gate_db_cnt_reg ( .CLK(clk), 
        .EN(N13), .ENCLK(net10992), .TE(1'b0) );
  DFFRQX1 db_cnt_reg_2_ ( .D(N16), .C(net10992), .XR(rstz), .Q(db_cnt[2]) );
  DFFRQX1 db_cnt_reg_1_ ( .D(N15), .C(net10992), .XR(rstz), .Q(db_cnt[1]) );
  DFFRQX1 db_cnt_reg_0_ ( .D(N14), .C(net10992), .XR(rstz), .Q(db_cnt[0]) );
  DFFRQX1 d_org_reg_0_ ( .D(i_org), .C(clk), .XR(rstz), .Q(d_org_0_) );
  DFFRQX1 d_org_reg_1_ ( .D(n7), .C(net10992), .XR(rstz), .Q(o_dbc) );
  OAI22X1 U3 ( .A(n4), .B(n1), .C(n6), .D(n3), .Y(N16) );
  INVX1 U4 ( .A(N14), .Y(n1) );
  NAND4X1 U5 ( .A(n5), .B(n2), .C(n3), .D(n4), .Y(N13) );
  XNOR2XL U6 ( .A(o_dbc), .B(d_org_0_), .Y(n5) );
  NOR4XL U7 ( .A(n4), .B(n2), .C(n5), .D(db_cnt[1]), .Y(o_chg) );
  INVX1 U8 ( .A(db_cnt[2]), .Y(n4) );
  INVX1 U9 ( .A(db_cnt[0]), .Y(n2) );
  AO22AXL U10 ( .A(d_org_0_), .B(o_chg), .C(o_dbc), .D(o_chg), .Y(n7) );
  NAND31X1 U11 ( .C(n5), .A(n4), .B(db_cnt[0]), .Y(n6) );
  NOR2X1 U12 ( .A(n5), .B(db_cnt[0]), .Y(N14) );
  OAI22X1 U13 ( .A(n3), .B(n1), .C(db_cnt[1]), .D(n6), .Y(N15) );
  INVX1 U14 ( .A(db_cnt[1]), .Y(n3) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dbnc_WIDTH3_TIMEOUT5_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module dbnc_WIDTH3_TIMEOUT5_2 ( o_dbc, o_chg, i_org, clk, rstz );
  input i_org, clk, rstz;
  output o_dbc, o_chg;
  wire   d_org_0_, N13, N14, N15, N16, net11010, n5, n6, n7, n1, n2, n3, n4;
  wire   [2:0] db_cnt;

  SNPS_CLOCK_GATE_HIGH_dbnc_WIDTH3_TIMEOUT5_2 clk_gate_db_cnt_reg ( .CLK(clk), 
        .EN(N13), .ENCLK(net11010), .TE(1'b0) );
  DFFRQX1 db_cnt_reg_2_ ( .D(N16), .C(net11010), .XR(rstz), .Q(db_cnt[2]) );
  DFFRQX1 db_cnt_reg_1_ ( .D(N15), .C(net11010), .XR(rstz), .Q(db_cnt[1]) );
  DFFRQX1 db_cnt_reg_0_ ( .D(N14), .C(net11010), .XR(rstz), .Q(db_cnt[0]) );
  DFFRQX1 d_org_reg_0_ ( .D(i_org), .C(clk), .XR(rstz), .Q(d_org_0_) );
  DFFRQX1 d_org_reg_1_ ( .D(n7), .C(net11010), .XR(rstz), .Q(o_dbc) );
  NOR4XL U3 ( .A(n4), .B(n2), .C(n5), .D(db_cnt[1]), .Y(o_chg) );
  OAI22X1 U4 ( .A(n4), .B(n1), .C(n6), .D(n3), .Y(N16) );
  INVX1 U5 ( .A(N14), .Y(n1) );
  NAND4X1 U6 ( .A(n5), .B(n2), .C(n3), .D(n4), .Y(N13) );
  XNOR2XL U7 ( .A(o_dbc), .B(d_org_0_), .Y(n5) );
  AO22AXL U8 ( .A(d_org_0_), .B(o_chg), .C(o_dbc), .D(o_chg), .Y(n7) );
  INVX1 U9 ( .A(db_cnt[2]), .Y(n4) );
  INVX1 U10 ( .A(db_cnt[0]), .Y(n2) );
  NAND31X1 U11 ( .C(n5), .A(n4), .B(db_cnt[0]), .Y(n6) );
  NOR2X1 U12 ( .A(n5), .B(db_cnt[0]), .Y(N14) );
  OAI22X1 U13 ( .A(n3), .B(n1), .C(db_cnt[1]), .D(n6), .Y(N15) );
  INVX1 U14 ( .A(db_cnt[1]), .Y(n3) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dbnc_WIDTH3_TIMEOUT5_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module dbnc_WIDTH3_TIMEOUT5_3 ( o_dbc, o_chg, i_org, clk, rstz );
  input i_org, clk, rstz;
  output o_dbc, o_chg;
  wire   d_org_0_, N13, N14, N15, N16, net11028, n5, n6, n7, n1, n2, n3, n4;
  wire   [2:0] db_cnt;

  SNPS_CLOCK_GATE_HIGH_dbnc_WIDTH3_TIMEOUT5_3 clk_gate_db_cnt_reg ( .CLK(clk), 
        .EN(N13), .ENCLK(net11028), .TE(1'b0) );
  DFFRQX1 db_cnt_reg_2_ ( .D(N16), .C(net11028), .XR(rstz), .Q(db_cnt[2]) );
  DFFRQX1 db_cnt_reg_1_ ( .D(N15), .C(net11028), .XR(rstz), .Q(db_cnt[1]) );
  DFFRQX1 d_org_reg_0_ ( .D(i_org), .C(clk), .XR(rstz), .Q(d_org_0_) );
  DFFRQX1 db_cnt_reg_0_ ( .D(N14), .C(net11028), .XR(rstz), .Q(db_cnt[0]) );
  DFFRQX1 d_org_reg_1_ ( .D(n7), .C(net11028), .XR(rstz), .Q(o_dbc) );
  NOR4XL U3 ( .A(n4), .B(n2), .C(n5), .D(db_cnt[1]), .Y(o_chg) );
  OAI22X1 U4 ( .A(n4), .B(n1), .C(n6), .D(n3), .Y(N16) );
  INVX1 U5 ( .A(N14), .Y(n1) );
  NAND4X1 U6 ( .A(n5), .B(n2), .C(n3), .D(n4), .Y(N13) );
  XNOR2XL U7 ( .A(o_dbc), .B(d_org_0_), .Y(n5) );
  INVX1 U8 ( .A(db_cnt[0]), .Y(n2) );
  AO22AXL U9 ( .A(d_org_0_), .B(o_chg), .C(o_dbc), .D(o_chg), .Y(n7) );
  INVX1 U10 ( .A(db_cnt[2]), .Y(n4) );
  NAND31X1 U11 ( .C(n5), .A(n4), .B(db_cnt[0]), .Y(n6) );
  NOR2X1 U12 ( .A(n5), .B(db_cnt[0]), .Y(N14) );
  OAI22X1 U13 ( .A(n3), .B(n1), .C(db_cnt[1]), .D(n6), .Y(N15) );
  INVX1 U14 ( .A(db_cnt[1]), .Y(n3) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dbnc_WIDTH3_TIMEOUT5_3 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module dbnc_WIDTH3_TIMEOUT5_4 ( o_dbc, o_chg, i_org, clk, rstz );
  input i_org, clk, rstz;
  output o_dbc, o_chg;
  wire   d_org_0_, N13, N14, N15, N16, net11046, n5, n6, n7, n1, n2, n3, n4;
  wire   [2:0] db_cnt;

  SNPS_CLOCK_GATE_HIGH_dbnc_WIDTH3_TIMEOUT5_4 clk_gate_db_cnt_reg ( .CLK(clk), 
        .EN(N13), .ENCLK(net11046), .TE(1'b0) );
  DFFRQX1 db_cnt_reg_2_ ( .D(N16), .C(net11046), .XR(rstz), .Q(db_cnt[2]) );
  DFFRQX1 db_cnt_reg_1_ ( .D(N15), .C(net11046), .XR(rstz), .Q(db_cnt[1]) );
  DFFRQX1 d_org_reg_0_ ( .D(i_org), .C(clk), .XR(rstz), .Q(d_org_0_) );
  DFFRQX1 db_cnt_reg_0_ ( .D(N14), .C(net11046), .XR(rstz), .Q(db_cnt[0]) );
  DFFRQX1 d_org_reg_1_ ( .D(n7), .C(net11046), .XR(rstz), .Q(o_dbc) );
  OAI22X1 U3 ( .A(n4), .B(n1), .C(n6), .D(n3), .Y(N16) );
  INVX1 U4 ( .A(N14), .Y(n1) );
  NAND4X1 U5 ( .A(n5), .B(n2), .C(n3), .D(n4), .Y(N13) );
  XNOR2XL U6 ( .A(o_dbc), .B(d_org_0_), .Y(n5) );
  NOR4XL U7 ( .A(n4), .B(n2), .C(n5), .D(db_cnt[1]), .Y(o_chg) );
  INVX1 U8 ( .A(db_cnt[0]), .Y(n2) );
  AO22AXL U9 ( .A(d_org_0_), .B(o_chg), .C(o_dbc), .D(o_chg), .Y(n7) );
  INVX1 U10 ( .A(db_cnt[2]), .Y(n4) );
  NAND31X1 U11 ( .C(n5), .A(n4), .B(db_cnt[0]), .Y(n6) );
  NOR2X1 U12 ( .A(n5), .B(db_cnt[0]), .Y(N14) );
  OAI22X1 U13 ( .A(n3), .B(n1), .C(db_cnt[1]), .D(n6), .Y(N15) );
  INVX1 U14 ( .A(db_cnt[1]), .Y(n3) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dbnc_WIDTH3_TIMEOUT5_4 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module dbnc_a0_2 ( o_dbc, o_chg, i_org, clk, rstz );
  input i_org, clk, rstz;
  output o_dbc, o_chg;
  wire   d_org_0_, N16, N17, N18, N19, N20, net11064, n5, n6, n7, n8, n9, n10,
         n11, n12, n1, n2, n3, n4;
  wire   [3:0] db_cnt;

  SNPS_CLOCK_GATE_HIGH_dbnc_a0_2 clk_gate_db_cnt_reg ( .CLK(clk), .EN(N16), 
        .ENCLK(net11064), .TE(1'b0) );
  DFFRQX1 d_org_reg_0_ ( .D(i_org), .C(clk), .XR(rstz), .Q(d_org_0_) );
  DFFRQX1 db_cnt_reg_3_ ( .D(N20), .C(net11064), .XR(rstz), .Q(db_cnt[3]) );
  DFFRQX1 db_cnt_reg_2_ ( .D(N19), .C(net11064), .XR(rstz), .Q(db_cnt[2]) );
  DFFRQX1 db_cnt_reg_1_ ( .D(N18), .C(net11064), .XR(rstz), .Q(db_cnt[1]) );
  DFFRQX1 db_cnt_reg_0_ ( .D(N17), .C(net11064), .XR(rstz), .Q(db_cnt[0]) );
  DFFRQX1 d_org_reg_1_ ( .D(n12), .C(net11064), .XR(rstz), .Q(o_dbc) );
  INVX1 U3 ( .A(n8), .Y(n1) );
  NOR21XL U4 ( .B(n5), .A(n6), .Y(o_chg) );
  NOR2X1 U5 ( .A(n3), .B(n7), .Y(n5) );
  NOR2X1 U6 ( .A(n6), .B(n5), .Y(n8) );
  OAI22X1 U7 ( .A(n1), .B(n3), .C(n7), .D(n1), .Y(N20) );
  NOR2X1 U8 ( .A(n10), .B(n1), .Y(N18) );
  XNOR2XL U9 ( .A(n4), .B(n2), .Y(n10) );
  NAND3X1 U10 ( .A(db_cnt[1]), .B(db_cnt[0]), .C(db_cnt[2]), .Y(n7) );
  XNOR2XL U11 ( .A(o_dbc), .B(d_org_0_), .Y(n6) );
  INVX1 U12 ( .A(db_cnt[3]), .Y(n3) );
  GEN2XL U13 ( .D(n8), .E(n4), .C(N17), .B(db_cnt[2]), .A(n9), .Y(N19) );
  NOR4XL U14 ( .A(db_cnt[2]), .B(n2), .C(n4), .D(n1), .Y(n9) );
  NOR2X1 U15 ( .A(n1), .B(db_cnt[0]), .Y(N17) );
  AO22AXL U16 ( .A(d_org_0_), .B(o_chg), .C(o_dbc), .D(o_chg), .Y(n12) );
  INVX1 U17 ( .A(db_cnt[0]), .Y(n2) );
  INVX1 U18 ( .A(db_cnt[1]), .Y(n4) );
  NAND3X1 U19 ( .A(n6), .B(n2), .C(n11), .Y(N16) );
  NOR3XL U20 ( .A(db_cnt[1]), .B(db_cnt[3]), .C(db_cnt[2]), .Y(n11) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dbnc_a0_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module dbnc_WIDTH4_TIMEOUT14_0 ( o_dbc, o_chg, i_org, clk, rstz );
  input i_org, clk, rstz;
  output o_dbc, o_chg;
  wire   d_org_0_, N15, N16, N17, N18, N19, net11082, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n1, n2, n3;
  wire   [3:0] db_cnt;

  SNPS_CLOCK_GATE_HIGH_dbnc_WIDTH4_TIMEOUT14_0 clk_gate_db_cnt_reg ( .CLK(clk), 
        .EN(N15), .ENCLK(net11082), .TE(1'b0) );
  DFFRQX1 db_cnt_reg_3_ ( .D(N19), .C(net11082), .XR(rstz), .Q(db_cnt[3]) );
  DFFRQX1 db_cnt_reg_0_ ( .D(N16), .C(net11082), .XR(rstz), .Q(db_cnt[0]) );
  DFFRQX1 d_org_reg_0_ ( .D(i_org), .C(clk), .XR(rstz), .Q(d_org_0_) );
  DFFRQX1 db_cnt_reg_1_ ( .D(N17), .C(net11082), .XR(rstz), .Q(db_cnt[1]) );
  DFFRQX1 db_cnt_reg_2_ ( .D(N18), .C(net11082), .XR(rstz), .Q(db_cnt[2]) );
  DFFRQX1 d_org_reg_1_ ( .D(n13), .C(net11082), .XR(rstz), .Q(o_dbc) );
  NAND21X1 U3 ( .B(n5), .A(n4), .Y(n7) );
  AOI21BBXL U4 ( .B(db_cnt[1]), .C(n7), .A(N16), .Y(n9) );
  XNOR2XL U5 ( .A(o_dbc), .B(d_org_0_), .Y(n5) );
  OAI32X1 U6 ( .A(n6), .B(n7), .C(n1), .D(n8), .E(n3), .Y(N19) );
  NAND3X1 U7 ( .A(db_cnt[1]), .B(n3), .C(db_cnt[2]), .Y(n6) );
  OA21X1 U8 ( .B(n7), .C(db_cnt[2]), .A(n9), .Y(n8) );
  INVX1 U9 ( .A(db_cnt[3]), .Y(n3) );
  NAND4X1 U10 ( .A(db_cnt[3]), .B(db_cnt[2]), .C(db_cnt[1]), .D(n1), .Y(n4) );
  NOR2X1 U11 ( .A(n7), .B(db_cnt[0]), .Y(N16) );
  AO22AXL U12 ( .A(d_org_0_), .B(o_chg), .C(o_dbc), .D(o_chg), .Y(n13) );
  NOR2X1 U13 ( .A(n4), .B(n5), .Y(o_chg) );
  OAI21X1 U14 ( .B(n9), .C(n2), .A(n10), .Y(N18) );
  NAND42X1 U15 ( .C(n7), .D(n1), .A(db_cnt[1]), .B(n2), .Y(n10) );
  INVX1 U16 ( .A(db_cnt[2]), .Y(n2) );
  INVX1 U17 ( .A(db_cnt[0]), .Y(n1) );
  NOR2X1 U18 ( .A(n11), .B(n7), .Y(N17) );
  XNOR2XL U19 ( .A(db_cnt[1]), .B(db_cnt[0]), .Y(n11) );
  NAND3X1 U20 ( .A(n5), .B(n1), .C(n12), .Y(N15) );
  NOR3XL U21 ( .A(db_cnt[1]), .B(db_cnt[3]), .C(db_cnt[2]), .Y(n12) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dbnc_WIDTH4_TIMEOUT14_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module dbnc_WIDTH4_TIMEOUT14_1 ( o_dbc, o_chg, i_org, clk, rstz );
  input i_org, clk, rstz;
  output o_dbc, o_chg;
  wire   d_org_0_, N15, N16, N17, N18, N19, net11100, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n1, n2, n3;
  wire   [3:0] db_cnt;

  SNPS_CLOCK_GATE_HIGH_dbnc_WIDTH4_TIMEOUT14_1 clk_gate_db_cnt_reg ( .CLK(clk), 
        .EN(N15), .ENCLK(net11100), .TE(1'b0) );
  DFFRQX1 db_cnt_reg_3_ ( .D(N19), .C(net11100), .XR(rstz), .Q(db_cnt[3]) );
  DFFRQX1 db_cnt_reg_0_ ( .D(N16), .C(net11100), .XR(rstz), .Q(db_cnt[0]) );
  DFFRQX1 d_org_reg_0_ ( .D(i_org), .C(clk), .XR(rstz), .Q(d_org_0_) );
  DFFRQX1 db_cnt_reg_1_ ( .D(N17), .C(net11100), .XR(rstz), .Q(db_cnt[1]) );
  DFFRQX1 db_cnt_reg_2_ ( .D(N18), .C(net11100), .XR(rstz), .Q(db_cnt[2]) );
  DFFRQX1 d_org_reg_1_ ( .D(n13), .C(net11100), .XR(rstz), .Q(o_dbc) );
  NAND21X1 U3 ( .B(n5), .A(n4), .Y(n7) );
  AOI21BBXL U4 ( .B(db_cnt[1]), .C(n7), .A(N16), .Y(n9) );
  XNOR2XL U5 ( .A(o_dbc), .B(d_org_0_), .Y(n5) );
  OAI32X1 U6 ( .A(n6), .B(n7), .C(n1), .D(n8), .E(n3), .Y(N19) );
  NAND3X1 U7 ( .A(db_cnt[1]), .B(n3), .C(db_cnt[2]), .Y(n6) );
  OA21X1 U8 ( .B(n7), .C(db_cnt[2]), .A(n9), .Y(n8) );
  INVX1 U9 ( .A(db_cnt[3]), .Y(n3) );
  NAND4X1 U10 ( .A(db_cnt[3]), .B(db_cnt[2]), .C(db_cnt[1]), .D(n1), .Y(n4) );
  NOR2X1 U11 ( .A(n7), .B(db_cnt[0]), .Y(N16) );
  AO22AXL U12 ( .A(d_org_0_), .B(o_chg), .C(o_dbc), .D(o_chg), .Y(n13) );
  NOR2X1 U13 ( .A(n4), .B(n5), .Y(o_chg) );
  OAI21X1 U14 ( .B(n9), .C(n2), .A(n10), .Y(N18) );
  NAND42X1 U15 ( .C(n7), .D(n1), .A(db_cnt[1]), .B(n2), .Y(n10) );
  INVX1 U16 ( .A(db_cnt[2]), .Y(n2) );
  INVX1 U17 ( .A(db_cnt[0]), .Y(n1) );
  NOR2X1 U18 ( .A(n11), .B(n7), .Y(N17) );
  XNOR2XL U19 ( .A(db_cnt[1]), .B(db_cnt[0]), .Y(n11) );
  NAND3X1 U20 ( .A(n5), .B(n1), .C(n12), .Y(N15) );
  NOR3XL U21 ( .A(db_cnt[1]), .B(db_cnt[3]), .C(db_cnt[2]), .Y(n12) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dbnc_WIDTH4_TIMEOUT14_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module dbnc_WIDTH4_TIMEOUT14_2 ( o_dbc, o_chg, i_org, clk, rstz );
  input i_org, clk, rstz;
  output o_dbc, o_chg;
  wire   d_org_0_, N15, N16, N17, N18, N19, net11118, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n1, n2, n3;
  wire   [3:0] db_cnt;

  SNPS_CLOCK_GATE_HIGH_dbnc_WIDTH4_TIMEOUT14_2 clk_gate_db_cnt_reg ( .CLK(clk), 
        .EN(N15), .ENCLK(net11118), .TE(1'b0) );
  DFFRQX1 db_cnt_reg_3_ ( .D(N19), .C(net11118), .XR(rstz), .Q(db_cnt[3]) );
  DFFRQX1 db_cnt_reg_0_ ( .D(N16), .C(net11118), .XR(rstz), .Q(db_cnt[0]) );
  DFFRQX1 d_org_reg_0_ ( .D(i_org), .C(clk), .XR(rstz), .Q(d_org_0_) );
  DFFRQX1 db_cnt_reg_1_ ( .D(N17), .C(net11118), .XR(rstz), .Q(db_cnt[1]) );
  DFFRQX1 db_cnt_reg_2_ ( .D(N18), .C(net11118), .XR(rstz), .Q(db_cnt[2]) );
  DFFRQX1 d_org_reg_1_ ( .D(n13), .C(net11118), .XR(rstz), .Q(o_dbc) );
  NAND21X1 U3 ( .B(n5), .A(n4), .Y(n7) );
  AOI21BBXL U4 ( .B(db_cnt[1]), .C(n7), .A(N16), .Y(n9) );
  XNOR2XL U5 ( .A(o_dbc), .B(d_org_0_), .Y(n5) );
  OAI32X1 U6 ( .A(n6), .B(n7), .C(n1), .D(n8), .E(n3), .Y(N19) );
  NAND3X1 U7 ( .A(db_cnt[1]), .B(n3), .C(db_cnt[2]), .Y(n6) );
  OA21X1 U8 ( .B(n7), .C(db_cnt[2]), .A(n9), .Y(n8) );
  INVX1 U9 ( .A(db_cnt[3]), .Y(n3) );
  NAND4X1 U10 ( .A(db_cnt[3]), .B(db_cnt[2]), .C(db_cnt[1]), .D(n1), .Y(n4) );
  NOR2X1 U11 ( .A(n7), .B(db_cnt[0]), .Y(N16) );
  AO22AXL U12 ( .A(d_org_0_), .B(o_chg), .C(o_dbc), .D(o_chg), .Y(n13) );
  NOR2X1 U13 ( .A(n4), .B(n5), .Y(o_chg) );
  OAI21X1 U14 ( .B(n9), .C(n2), .A(n10), .Y(N18) );
  NAND42X1 U15 ( .C(n7), .D(n1), .A(db_cnt[1]), .B(n2), .Y(n10) );
  INVX1 U16 ( .A(db_cnt[2]), .Y(n2) );
  INVX1 U17 ( .A(db_cnt[0]), .Y(n1) );
  NOR2X1 U18 ( .A(n11), .B(n7), .Y(N17) );
  XNOR2XL U19 ( .A(db_cnt[1]), .B(db_cnt[0]), .Y(n11) );
  NAND3X1 U20 ( .A(n5), .B(n1), .C(n12), .Y(N15) );
  NOR3XL U21 ( .A(db_cnt[1]), .B(db_cnt[3]), .C(db_cnt[2]), .Y(n12) );
endmodule


module SNPS_CLOCK_GATE_HIGH_dbnc_WIDTH4_TIMEOUT14_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_8_00000028 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net11136;

  SNPS_CLOCK_GATE_HIGH_glreg_8_00000028 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11136), .TE(1'b0) );
  DFFSQX1 mem_reg_5_ ( .D(wdat[5]), .C(net11136), .XS(arstz), .Q(rdat[5]) );
  DFFSQX1 mem_reg_3_ ( .D(wdat[3]), .C(net11136), .XS(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net11136), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net11136), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net11136), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net11136), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net11136), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net11136), .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_8_00000028 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_56 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net11154;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_56 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11154), .TE(1'b0) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net11154), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net11154), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net11154), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net11154), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net11154), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net11154), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net11154), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net11154), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_56 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_57 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net11172;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_57 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11172), .TE(1'b0) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net11172), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net11172), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net11172), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net11172), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net11172), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net11172), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net11172), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net11172), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_57 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_58 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net11190;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_58 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11190), .TE(1'b0) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net11190), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net11190), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net11190), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net11190), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net11190), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net11190), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net11190), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net11190), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_58 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_59 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net11208;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_59 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11208), .TE(1'b0) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net11208), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net11208), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net11208), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net11208), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net11208), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net11208), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net11208), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net11208), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_59 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_60 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net11226;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_60 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11226), .TE(1'b0) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net11226), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net11226), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net11226), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net11226), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net11226), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net11226), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net11226), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net11226), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_60 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_61 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net11244;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_61 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11244), .TE(1'b0) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net11244), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net11244), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net11244), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net11244), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net11244), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net11244), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net11244), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net11244), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_61 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_62 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net11262;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_62 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11262), .TE(1'b0) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net11262), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net11262), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net11262), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net11262), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net11262), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net11262), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net11262), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net11262), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_62 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_63 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net11280;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_63 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11280), .TE(1'b0) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net11280), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net11280), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net11280), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net11280), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net11280), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net11280), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net11280), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net11280), .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_63 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_WIDTH4 ( clk, arstz, we, wdat, rdat );
  input [3:0] wdat;
  output [3:0] rdat;
  input clk, arstz, we;
  wire   net11298;

  SNPS_CLOCK_GATE_HIGH_glreg_WIDTH4 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11298), .TE(1'b0) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net11298), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net11298), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net11298), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net11298), .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_WIDTH4 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_64 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net11316;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_64 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11316), .TE(1'b0) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net11316), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net11316), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net11316), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net11316), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net11316), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net11316), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net11316), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net11316), .XR(arstz), .Q(rdat[2]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_64 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glsta_a0_3 ( clk, arstz, rst0, set2, clr1, rdat, irq );
  input [7:0] set2;
  input [7:0] clr1;
  output [7:0] rdat;
  output [7:0] irq;
  input clk, arstz, rst0;
  wire   upd_r, n17, n18, n19, n20, n21, n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16;
  wire   [7:0] wd_r;

  glreg_WIDTH8_3 u0 ( .clk(clk), .arstz(arstz), .we(upd_r), .wdat(wd_r), 
        .rdat(rdat) );
  NOR4XL U2 ( .A(clr1[7]), .B(clr1[6]), .C(clr1[5]), .D(clr1[4]), .Y(n18) );
  INVX1 U3 ( .A(set2[0]), .Y(n16) );
  INVX1 U4 ( .A(set2[1]), .Y(n15) );
  INVX1 U5 ( .A(set2[2]), .Y(n14) );
  INVX1 U6 ( .A(set2[3]), .Y(n13) );
  INVX1 U7 ( .A(set2[4]), .Y(n12) );
  NAND3X1 U8 ( .A(n10), .B(n9), .C(n11), .Y(n21) );
  NAND4X1 U9 ( .A(n17), .B(n18), .C(n19), .D(n20), .Y(upd_r) );
  NOR4XL U10 ( .A(set2[2]), .B(set2[1]), .C(set2[0]), .D(rst0), .Y(n19) );
  NOR3XL U11 ( .A(n21), .B(set2[4]), .C(set2[3]), .Y(n20) );
  NOR4XL U12 ( .A(clr1[3]), .B(clr1[2]), .C(clr1[1]), .D(clr1[0]), .Y(n17) );
  AOI211X1 U13 ( .C(n16), .D(n8), .A(rst0), .B(clr1[0]), .Y(wd_r[0]) );
  INVX1 U14 ( .A(rdat[0]), .Y(n8) );
  AOI211X1 U15 ( .C(n15), .D(n7), .A(rst0), .B(clr1[1]), .Y(wd_r[1]) );
  INVX1 U16 ( .A(rdat[1]), .Y(n7) );
  AOI211X1 U17 ( .C(n14), .D(n6), .A(rst0), .B(clr1[2]), .Y(wd_r[2]) );
  INVX1 U18 ( .A(rdat[2]), .Y(n6) );
  AOI211X1 U19 ( .C(n13), .D(n5), .A(rst0), .B(clr1[3]), .Y(wd_r[3]) );
  INVX1 U20 ( .A(rdat[3]), .Y(n5) );
  AOI211X1 U21 ( .C(n12), .D(n4), .A(rst0), .B(clr1[4]), .Y(wd_r[4]) );
  INVX1 U22 ( .A(rdat[4]), .Y(n4) );
  AOI211X1 U23 ( .C(n11), .D(n3), .A(rst0), .B(clr1[5]), .Y(wd_r[5]) );
  INVX1 U24 ( .A(rdat[5]), .Y(n3) );
  AOI211X1 U25 ( .C(n10), .D(n2), .A(rst0), .B(clr1[6]), .Y(wd_r[6]) );
  INVX1 U26 ( .A(rdat[6]), .Y(n2) );
  AOI211X1 U27 ( .C(n9), .D(n1), .A(rst0), .B(clr1[7]), .Y(wd_r[7]) );
  INVX1 U28 ( .A(rdat[7]), .Y(n1) );
  NOR2X1 U29 ( .A(rdat[0]), .B(n16), .Y(irq[0]) );
  NOR2X1 U30 ( .A(rdat[1]), .B(n15), .Y(irq[1]) );
  NOR2X1 U31 ( .A(rdat[2]), .B(n14), .Y(irq[2]) );
  NOR2X1 U32 ( .A(rdat[3]), .B(n13), .Y(irq[3]) );
  INVX1 U33 ( .A(set2[6]), .Y(n10) );
  INVX1 U34 ( .A(set2[7]), .Y(n9) );
  INVX1 U35 ( .A(set2[5]), .Y(n11) );
  NOR2X1 U36 ( .A(rdat[4]), .B(n12), .Y(irq[4]) );
  NOR2X1 U37 ( .A(rdat[6]), .B(n10), .Y(irq[6]) );
  NOR2X1 U38 ( .A(rdat[5]), .B(n11), .Y(irq[5]) );
  NOR2X1 U39 ( .A(rdat[7]), .B(n9), .Y(irq[7]) );
endmodule


module glreg_WIDTH8_3 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net11334;

  SNPS_CLOCK_GATE_HIGH_glreg_WIDTH8_3 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11334), .TE(1'b0) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net11334), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net11334), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net11334), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net11334), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net11334), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net11334), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net11334), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net11334), .XR(arstz), .Q(rdat[4]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_WIDTH8_3 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_65 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net11352;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_65 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11352), .TE(1'b0) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net11352), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net11352), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net11352), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net11352), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net11352), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net11352), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net11352), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net11352), .XR(arstz), .Q(rdat[4]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_65 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_66 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net11370;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_66 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11370), .TE(1'b0) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net11370), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net11370), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net11370), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net11370), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net11370), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net11370), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net11370), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net11370), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_66 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_8_00000032 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net11388;

  SNPS_CLOCK_GATE_HIGH_glreg_8_00000032 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11388), .TE(1'b0) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net11388), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net11388), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net11388), .XR(arstz), .Q(rdat[2]) );
  DFFSQX1 mem_reg_5_ ( .D(wdat[5]), .C(net11388), .XS(arstz), .Q(rdat[5]) );
  DFFSQX1 mem_reg_1_ ( .D(wdat[1]), .C(net11388), .XS(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net11388), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net11388), .XR(arstz), .Q(rdat[0]) );
  DFFSQX1 mem_reg_4_ ( .D(wdat[4]), .C(net11388), .XS(arstz), .Q(rdat[4]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_8_00000032 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_8_00000098 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net11406;

  SNPS_CLOCK_GATE_HIGH_glreg_8_00000098 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11406), .TE(1'b0) );
  DFFSQX1 mem_reg_7_ ( .D(wdat[7]), .C(net11406), .XS(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net11406), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net11406), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net11406), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net11406), .XR(arstz), .Q(rdat[0]) );
  DFFSQX1 mem_reg_3_ ( .D(wdat[3]), .C(net11406), .XS(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net11406), .XR(arstz), .Q(rdat[1]) );
  DFFSQX1 mem_reg_4_ ( .D(wdat[4]), .C(net11406), .XS(arstz), .Q(rdat[4]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_8_00000098 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_8_000000f0 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net11424;

  SNPS_CLOCK_GATE_HIGH_glreg_8_000000f0 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11424), .TE(1'b0) );
  DFFSQX1 mem_reg_7_ ( .D(wdat[7]), .C(net11424), .XS(arstz), .Q(rdat[7]) );
  DFFSQX1 mem_reg_6_ ( .D(wdat[6]), .C(net11424), .XS(arstz), .Q(rdat[6]) );
  DFFSQX1 mem_reg_5_ ( .D(wdat[5]), .C(net11424), .XS(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net11424), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net11424), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net11424), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net11424), .XR(arstz), .Q(rdat[0]) );
  DFFSQX1 mem_reg_4_ ( .D(wdat[4]), .C(net11424), .XS(arstz), .Q(rdat[4]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_8_000000f0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_WIDTH1_3 ( clk, arstz, we, wdat, rdat );
  input [0:0] wdat;
  output [0:0] rdat;
  input clk, arstz, we;
  wire   n2;

  DFFRQX1 mem_reg_0_ ( .D(n2), .C(clk), .XR(arstz), .Q(rdat[0]) );
  AO22AXL U2 ( .A(we), .B(wdat[0]), .C(rdat[0]), .D(we), .Y(n2) );
endmodule


module glreg_WIDTH1_4 ( clk, arstz, we, wdat, rdat );
  input [0:0] wdat;
  output [0:0] rdat;
  input clk, arstz, we;
  wire   n2;

  DFFRQX1 mem_reg_0_ ( .D(n2), .C(clk), .XR(arstz), .Q(rdat[0]) );
  AO22AXL U2 ( .A(we), .B(wdat[0]), .C(rdat[0]), .D(we), .Y(n2) );
endmodule


module glreg_WIDTH1_5 ( clk, arstz, we, wdat, rdat );
  input [0:0] wdat;
  output [0:0] rdat;
  input clk, arstz, we;
  wire   n2;

  DFFRQX1 mem_reg_0_ ( .D(n2), .C(clk), .XR(arstz), .Q(rdat[0]) );
  AO22AXL U2 ( .A(we), .B(wdat[0]), .C(rdat[0]), .D(we), .Y(n2) );
endmodule


module glreg_WIDTH2_2 ( clk, arstz, we, wdat, rdat );
  input [1:0] wdat;
  output [1:0] rdat;
  input clk, arstz, we;
  wire   n2, n3, n1;

  DFFRQX1 mem_reg_0_ ( .D(n2), .C(clk), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_1_ ( .D(n3), .C(clk), .XR(arstz), .Q(rdat[1]) );
  INVXL U2 ( .A(we), .Y(n1) );
  AO22XL U3 ( .A(we), .B(wdat[0]), .C(rdat[0]), .D(n1), .Y(n2) );
  AO22XL U4 ( .A(wdat[1]), .B(we), .C(rdat[1]), .D(n1), .Y(n3) );
endmodule


module glreg_WIDTH3 ( clk, arstz, we, wdat, rdat );
  input [2:0] wdat;
  output [2:0] rdat;
  input clk, arstz, we;
  wire   net11442;

  SNPS_CLOCK_GATE_HIGH_glreg_WIDTH3 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11442), .TE(1'b0) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net11442), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net11442), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net11442), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_WIDTH3 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_8_00000011 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net11460;

  SNPS_CLOCK_GATE_HIGH_glreg_8_00000011 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11460), .TE(1'b0) );
  DFFSQX1 mem_reg_4_ ( .D(wdat[4]), .C(net11460), .XS(arstz), .Q(rdat[4]) );
  DFFSQX1 mem_reg_0_ ( .D(wdat[0]), .C(net11460), .XS(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net11460), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net11460), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net11460), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net11460), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net11460), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net11460), .XR(arstz), .Q(rdat[3]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_8_00000011 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_8_00000001 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net11478;

  SNPS_CLOCK_GATE_HIGH_glreg_8_00000001 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11478), .TE(1'b0) );
  DFFSQX1 mem_reg_0_ ( .D(wdat[0]), .C(net11478), .XS(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net11478), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net11478), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net11478), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net11478), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net11478), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net11478), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net11478), .XR(arstz), .Q(rdat[6]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_8_00000001 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_67 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net11496;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_67 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11496), .TE(1'b0) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net11496), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net11496), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net11496), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net11496), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net11496), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net11496), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net11496), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net11496), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_67 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glsta_a0_4 ( clk, arstz, rst0, set2, clr1, rdat, irq );
  input [7:0] set2;
  input [7:0] clr1;
  output [7:0] rdat;
  output [7:0] irq;
  input clk, arstz, rst0;
  wire   upd_r, n17, n18, n19, n20, n21, n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16;
  wire   [7:0] wd_r;

  glreg_WIDTH8_4 u0 ( .clk(clk), .arstz(arstz), .we(upd_r), .wdat(wd_r), 
        .rdat(rdat) );
  NOR4XL U2 ( .A(clr1[7]), .B(clr1[6]), .C(clr1[5]), .D(clr1[4]), .Y(n18) );
  NAND3X1 U3 ( .A(n3), .B(n4), .C(n2), .Y(n21) );
  INVX1 U4 ( .A(set2[3]), .Y(n14) );
  INVX1 U5 ( .A(set2[1]), .Y(n16) );
  INVX1 U6 ( .A(set2[0]), .Y(n13) );
  INVX1 U7 ( .A(set2[4]), .Y(n1) );
  INVX1 U8 ( .A(set2[6]), .Y(n3) );
  INVX1 U9 ( .A(set2[7]), .Y(n4) );
  INVX1 U10 ( .A(set2[2]), .Y(n15) );
  INVX1 U11 ( .A(set2[5]), .Y(n2) );
  NAND4X1 U12 ( .A(n17), .B(n18), .C(n19), .D(n20), .Y(upd_r) );
  NOR4XL U13 ( .A(set2[2]), .B(set2[1]), .C(set2[0]), .D(rst0), .Y(n19) );
  NOR3XL U14 ( .A(n21), .B(set2[4]), .C(set2[3]), .Y(n20) );
  NOR4XL U15 ( .A(clr1[3]), .B(clr1[2]), .C(clr1[1]), .D(clr1[0]), .Y(n17) );
  AOI211X1 U16 ( .C(n13), .D(n12), .A(rst0), .B(clr1[0]), .Y(wd_r[0]) );
  INVX1 U17 ( .A(rdat[0]), .Y(n12) );
  AOI211X1 U18 ( .C(n16), .D(n11), .A(rst0), .B(clr1[1]), .Y(wd_r[1]) );
  INVX1 U19 ( .A(rdat[1]), .Y(n11) );
  AOI211X1 U20 ( .C(n15), .D(n10), .A(rst0), .B(clr1[2]), .Y(wd_r[2]) );
  INVX1 U21 ( .A(rdat[2]), .Y(n10) );
  AOI211X1 U22 ( .C(n14), .D(n9), .A(rst0), .B(clr1[3]), .Y(wd_r[3]) );
  INVX1 U23 ( .A(rdat[3]), .Y(n9) );
  AOI211X1 U24 ( .C(n1), .D(n8), .A(rst0), .B(clr1[4]), .Y(wd_r[4]) );
  INVX1 U25 ( .A(rdat[4]), .Y(n8) );
  AOI211X1 U26 ( .C(n2), .D(n7), .A(rst0), .B(clr1[5]), .Y(wd_r[5]) );
  INVX1 U27 ( .A(rdat[5]), .Y(n7) );
  AOI211X1 U28 ( .C(n3), .D(n6), .A(rst0), .B(clr1[6]), .Y(wd_r[6]) );
  INVX1 U29 ( .A(rdat[6]), .Y(n6) );
  AOI211X1 U30 ( .C(n4), .D(n5), .A(rst0), .B(clr1[7]), .Y(wd_r[7]) );
  INVX1 U31 ( .A(rdat[7]), .Y(n5) );
  NOR2X1 U32 ( .A(rdat[7]), .B(n4), .Y(irq[7]) );
  NOR2X1 U33 ( .A(rdat[6]), .B(n3), .Y(irq[6]) );
  NOR2X1 U34 ( .A(rdat[3]), .B(n14), .Y(irq[3]) );
  NOR2X1 U35 ( .A(rdat[2]), .B(n15), .Y(irq[2]) );
  NOR2X1 U36 ( .A(rdat[0]), .B(n13), .Y(irq[0]) );
  NOR2X1 U37 ( .A(rdat[4]), .B(n1), .Y(irq[4]) );
  NOR2X1 U38 ( .A(rdat[5]), .B(n2), .Y(irq[5]) );
  NOR2X1 U39 ( .A(rdat[1]), .B(n16), .Y(irq[1]) );
endmodule


module glreg_WIDTH8_4 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net11514;

  SNPS_CLOCK_GATE_HIGH_glreg_WIDTH8_4 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11514), .TE(1'b0) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net11514), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net11514), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net11514), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net11514), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net11514), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net11514), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net11514), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net11514), .XR(arstz), .Q(rdat[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_WIDTH8_4 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_68 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net11532;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_68 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11532), .TE(1'b0) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net11532), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net11532), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net11532), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net11532), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net11532), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net11532), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net11532), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net11532), .XR(arstz), .Q(rdat[6]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_68 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_7_70 ( clk, arstz, we, wdat, rdat );
  input [6:0] wdat;
  output [6:0] rdat;
  input clk, arstz, we;
  wire   net11550;

  SNPS_CLOCK_GATE_HIGH_glreg_7_70 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11550), .TE(1'b0) );
  DFFSQX1 mem_reg_4_ ( .D(wdat[4]), .C(net11550), .XS(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net11550), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net11550), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net11550), .XR(arstz), .Q(rdat[0]) );
  DFFSQX1 mem_reg_6_ ( .D(wdat[6]), .C(net11550), .XS(arstz), .Q(rdat[6]) );
  DFFSQX1 mem_reg_5_ ( .D(wdat[5]), .C(net11550), .XS(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net11550), .XR(arstz), .Q(rdat[3]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_7_70 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_1_1 ( clk, arstz, we, wdat, rdat );
  input [0:0] wdat;
  output [0:0] rdat;
  input clk, arstz, we;
  wire   n1;

  DFFSQX1 mem_reg_0_ ( .D(n1), .C(clk), .XS(arstz), .Q(rdat[0]) );
  AO22AXL U2 ( .A(we), .B(wdat[0]), .C(rdat[0]), .D(we), .Y(n1) );
endmodule


module glreg_WIDTH1_6 ( clk, arstz, we, wdat, rdat );
  input [0:0] wdat;
  output [0:0] rdat;
  input clk, arstz, we;
  wire   n1;

  DFFRQX1 mem_reg_0_ ( .D(n1), .C(clk), .XR(arstz), .Q(rdat[0]) );
  AO22AXL U2 ( .A(we), .B(wdat[0]), .C(rdat[0]), .D(we), .Y(n1) );
endmodule


module glreg_6_00000018 ( clk, arstz, we, wdat, rdat );
  input [5:0] wdat;
  output [5:0] rdat;
  input clk, arstz, we;
  wire   net11568;

  SNPS_CLOCK_GATE_HIGH_glreg_6_00000018 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11568), .TE(1'b0) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net11568), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net11568), .XR(arstz), .Q(rdat[5]) );
  DFFSQX1 mem_reg_4_ ( .D(wdat[4]), .C(net11568), .XS(arstz), .Q(rdat[4]) );
  DFFSQX1 mem_reg_3_ ( .D(wdat[3]), .C(net11568), .XS(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net11568), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net11568), .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_6_00000018 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_69 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net11586;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_69 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11586), .TE(1'b0) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net11586), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net11586), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net11586), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net11586), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net11586), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net11586), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net11586), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net11586), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_69 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_70 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net11604;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_70 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11604), .TE(1'b0) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net11604), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net11604), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net11604), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net11604), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net11604), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net11604), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net11604), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net11604), .XR(arstz), .Q(rdat[6]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_70 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_71 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net11622;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_71 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11622), .TE(1'b0) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net11622), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net11622), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net11622), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net11622), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net11622), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net11622), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net11622), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net11622), .XR(arstz), .Q(rdat[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_71 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_72 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net11640;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_72 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11640), .TE(1'b0) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net11640), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net11640), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net11640), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net11640), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net11640), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net11640), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net11640), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net11640), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_72 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_73 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net11658;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_73 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11658), .TE(1'b0) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net11658), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net11658), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net11658), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net11658), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net11658), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net11658), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net11658), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net11658), .XR(arstz), .Q(rdat[4]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_73 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_WIDTH5_2 ( clk, arstz, we, wdat, rdat );
  input [4:0] wdat;
  output [4:0] rdat;
  input clk, arstz, we;
  wire   net11676;

  SNPS_CLOCK_GATE_HIGH_glreg_WIDTH5_2 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11676), .TE(1'b0) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net11676), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net11676), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net11676), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net11676), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net11676), .XR(arstz), .Q(rdat[2]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_WIDTH5_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_74 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net11694;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_74 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11694), .TE(1'b0) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net11694), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net11694), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net11694), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net11694), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net11694), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net11694), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net11694), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net11694), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_74 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_75 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net11712;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_75 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11712), .TE(1'b0) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net11712), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net11712), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net11712), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net11712), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net11712), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net11712), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net11712), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net11712), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_75 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_76 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net11730;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_76 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11730), .TE(1'b0) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net11730), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net11730), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net11730), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net11730), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net11730), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net11730), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net11730), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net11730), .XR(arstz), .Q(rdat[4]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_76 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_77 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net11748;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_77 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11748), .TE(1'b0) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net11748), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net11748), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net11748), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net11748), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net11748), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net11748), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net11748), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net11748), .XR(arstz), .Q(rdat[4]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_77 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glsta_a0_5 ( clk, arstz, rst0, set2, clr1, rdat, irq );
  input [7:0] set2;
  input [7:0] clr1;
  output [7:0] rdat;
  output [7:0] irq;
  input clk, arstz, rst0;
  wire   upd_r, n17, n18, n19, n20, n21, n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16;
  wire   [7:0] wd_r;

  glreg_WIDTH8_5 u0 ( .clk(clk), .arstz(arstz), .we(upd_r), .wdat(wd_r), 
        .rdat(rdat) );
  NOR3XL U2 ( .A(n21), .B(set2[4]), .C(set2[3]), .Y(n20) );
  NAND3X1 U3 ( .A(n14), .B(n3), .C(n2), .Y(n21) );
  INVX1 U4 ( .A(set2[4]), .Y(n1) );
  INVX1 U5 ( .A(set2[3]), .Y(n4) );
  INVX1 U6 ( .A(set2[1]), .Y(n15) );
  INVX1 U7 ( .A(set2[2]), .Y(n5) );
  INVX1 U8 ( .A(set2[5]), .Y(n2) );
  NAND4X1 U9 ( .A(n17), .B(n18), .C(n19), .D(n20), .Y(upd_r) );
  NOR4XL U10 ( .A(clr1[3]), .B(clr1[2]), .C(clr1[1]), .D(clr1[0]), .Y(n17) );
  NOR4XL U11 ( .A(clr1[7]), .B(clr1[6]), .C(clr1[5]), .D(clr1[4]), .Y(n18) );
  NOR4XL U12 ( .A(set2[2]), .B(set2[1]), .C(set2[0]), .D(rst0), .Y(n19) );
  INVX1 U13 ( .A(set2[6]), .Y(n14) );
  INVX1 U14 ( .A(set2[0]), .Y(n16) );
  INVX1 U15 ( .A(set2[7]), .Y(n3) );
  NOR2X1 U16 ( .A(rdat[4]), .B(n1), .Y(irq[4]) );
  NOR2X1 U17 ( .A(rdat[5]), .B(n2), .Y(irq[5]) );
  AOI211X1 U18 ( .C(n1), .D(n9), .A(rst0), .B(clr1[4]), .Y(wd_r[4]) );
  INVX1 U19 ( .A(rdat[4]), .Y(n9) );
  AOI211X1 U20 ( .C(n2), .D(n8), .A(rst0), .B(clr1[5]), .Y(wd_r[5]) );
  INVX1 U21 ( .A(rdat[5]), .Y(n8) );
  AOI211X1 U22 ( .C(n16), .D(n13), .A(rst0), .B(clr1[0]), .Y(wd_r[0]) );
  INVX1 U23 ( .A(rdat[0]), .Y(n13) );
  AOI211X1 U24 ( .C(n15), .D(n12), .A(rst0), .B(clr1[1]), .Y(wd_r[1]) );
  INVX1 U25 ( .A(rdat[1]), .Y(n12) );
  AOI211X1 U26 ( .C(n5), .D(n11), .A(rst0), .B(clr1[2]), .Y(wd_r[2]) );
  INVX1 U27 ( .A(rdat[2]), .Y(n11) );
  AOI211X1 U28 ( .C(n4), .D(n10), .A(rst0), .B(clr1[3]), .Y(wd_r[3]) );
  INVX1 U29 ( .A(rdat[3]), .Y(n10) );
  AOI211X1 U30 ( .C(n14), .D(n7), .A(rst0), .B(clr1[6]), .Y(wd_r[6]) );
  INVX1 U31 ( .A(rdat[6]), .Y(n7) );
  AOI211X1 U32 ( .C(n3), .D(n6), .A(rst0), .B(clr1[7]), .Y(wd_r[7]) );
  INVX1 U33 ( .A(rdat[7]), .Y(n6) );
  NOR2X1 U34 ( .A(rdat[2]), .B(n5), .Y(irq[2]) );
  NOR2X1 U35 ( .A(rdat[3]), .B(n4), .Y(irq[3]) );
  NOR2X1 U36 ( .A(rdat[0]), .B(n16), .Y(irq[0]) );
  NOR2X1 U37 ( .A(rdat[6]), .B(n14), .Y(irq[6]) );
  NOR2X1 U38 ( .A(rdat[1]), .B(n15), .Y(irq[1]) );
  NOR2X1 U39 ( .A(rdat[7]), .B(n3), .Y(irq[7]) );
endmodule


module glreg_WIDTH8_5 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net11766;

  SNPS_CLOCK_GATE_HIGH_glreg_WIDTH8_5 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11766), .TE(1'b0) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net11766), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net11766), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net11766), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net11766), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net11766), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net11766), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net11766), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net11766), .XR(arstz), .Q(rdat[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_WIDTH8_5 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glsta_a0_6 ( clk, arstz, rst0, set2, clr1, rdat, irq );
  input [7:0] set2;
  input [7:0] clr1;
  output [7:0] rdat;
  output [7:0] irq;
  input clk, arstz, rst0;
  wire   upd_r, n17, n18, n19, n20, n21, n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16;
  wire   [7:0] wd_r;

  glreg_WIDTH8_6 u0 ( .clk(clk), .arstz(arstz), .we(upd_r), .wdat(wd_r), 
        .rdat(rdat) );
  INVX1 U2 ( .A(set2[7]), .Y(n2) );
  INVX1 U3 ( .A(set2[3]), .Y(n5) );
  INVX1 U4 ( .A(set2[1]), .Y(n1) );
  INVX1 U5 ( .A(set2[2]), .Y(n3) );
  INVX1 U6 ( .A(set2[4]), .Y(n6) );
  NOR3XL U7 ( .A(n21), .B(set2[4]), .C(set2[3]), .Y(n20) );
  NAND3X1 U8 ( .A(n4), .B(n2), .C(n15), .Y(n21) );
  NAND4X1 U9 ( .A(n17), .B(n18), .C(n19), .D(n20), .Y(upd_r) );
  NOR4XL U10 ( .A(clr1[3]), .B(clr1[2]), .C(clr1[1]), .D(clr1[0]), .Y(n17) );
  NOR4XL U11 ( .A(clr1[7]), .B(clr1[6]), .C(clr1[5]), .D(clr1[4]), .Y(n18) );
  NOR4XL U12 ( .A(set2[2]), .B(set2[1]), .C(set2[0]), .D(rst0), .Y(n19) );
  INVX1 U13 ( .A(set2[6]), .Y(n4) );
  INVX1 U14 ( .A(set2[0]), .Y(n16) );
  NOR2X1 U15 ( .A(rdat[6]), .B(n4), .Y(irq[6]) );
  NOR2X1 U16 ( .A(rdat[7]), .B(n2), .Y(irq[7]) );
  NOR2X1 U17 ( .A(rdat[2]), .B(n3), .Y(irq[2]) );
  NOR2X1 U18 ( .A(rdat[0]), .B(n16), .Y(irq[0]) );
  NOR2X1 U19 ( .A(rdat[1]), .B(n1), .Y(irq[1]) );
  AOI211X1 U20 ( .C(n2), .D(n7), .A(rst0), .B(clr1[7]), .Y(wd_r[7]) );
  INVX1 U21 ( .A(rdat[7]), .Y(n7) );
  AOI211X1 U22 ( .C(n16), .D(n14), .A(rst0), .B(clr1[0]), .Y(wd_r[0]) );
  INVX1 U23 ( .A(rdat[0]), .Y(n14) );
  AOI211X1 U24 ( .C(n4), .D(n8), .A(rst0), .B(clr1[6]), .Y(wd_r[6]) );
  INVX1 U25 ( .A(rdat[6]), .Y(n8) );
  AOI211X1 U26 ( .C(n1), .D(n13), .A(rst0), .B(clr1[1]), .Y(wd_r[1]) );
  INVX1 U27 ( .A(rdat[1]), .Y(n13) );
  AOI211X1 U28 ( .C(n3), .D(n12), .A(rst0), .B(clr1[2]), .Y(wd_r[2]) );
  INVX1 U29 ( .A(rdat[2]), .Y(n12) );
  AOI211X1 U30 ( .C(n5), .D(n11), .A(rst0), .B(clr1[3]), .Y(wd_r[3]) );
  INVX1 U31 ( .A(rdat[3]), .Y(n11) );
  AOI211X1 U32 ( .C(n6), .D(n10), .A(rst0), .B(clr1[4]), .Y(wd_r[4]) );
  INVX1 U33 ( .A(rdat[4]), .Y(n10) );
  AOI211X1 U34 ( .C(n15), .D(n9), .A(rst0), .B(clr1[5]), .Y(wd_r[5]) );
  INVX1 U35 ( .A(rdat[5]), .Y(n9) );
  NOR2X1 U36 ( .A(rdat[4]), .B(n6), .Y(irq[4]) );
  NOR2X1 U37 ( .A(rdat[3]), .B(n5), .Y(irq[3]) );
  INVX1 U38 ( .A(set2[5]), .Y(n15) );
  NOR2X1 U39 ( .A(rdat[5]), .B(n15), .Y(irq[5]) );
endmodule


module glreg_WIDTH8_6 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net11784;

  SNPS_CLOCK_GATE_HIGH_glreg_WIDTH8_6 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11784), .TE(1'b0) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net11784), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net11784), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net11784), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net11784), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net11784), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net11784), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net11784), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net11784), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_WIDTH8_6 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_78 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net11802;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_78 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11802), .TE(1'b0) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net11802), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net11802), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net11802), .XR(arstz), .Q(rdat[7]) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net11802), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net11802), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net11802), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net11802), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net11802), .XR(arstz), .Q(rdat[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_78 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module glreg_a0_79 ( clk, arstz, we, wdat, rdat );
  input [7:0] wdat;
  output [7:0] rdat;
  input clk, arstz, we;
  wire   net11820;

  SNPS_CLOCK_GATE_HIGH_glreg_a0_79 clk_gate_mem_reg ( .CLK(clk), .EN(we), 
        .ENCLK(net11820), .TE(1'b0) );
  DFFRQX1 mem_reg_4_ ( .D(wdat[4]), .C(net11820), .XR(arstz), .Q(rdat[4]) );
  DFFRQX1 mem_reg_2_ ( .D(wdat[2]), .C(net11820), .XR(arstz), .Q(rdat[2]) );
  DFFRQX1 mem_reg_1_ ( .D(wdat[1]), .C(net11820), .XR(arstz), .Q(rdat[1]) );
  DFFRQX1 mem_reg_0_ ( .D(wdat[0]), .C(net11820), .XR(arstz), .Q(rdat[0]) );
  DFFRQX1 mem_reg_5_ ( .D(wdat[5]), .C(net11820), .XR(arstz), .Q(rdat[5]) );
  DFFRQX1 mem_reg_3_ ( .D(wdat[3]), .C(net11820), .XR(arstz), .Q(rdat[3]) );
  DFFRQX1 mem_reg_6_ ( .D(wdat[6]), .C(net11820), .XR(arstz), .Q(rdat[6]) );
  DFFRQX1 mem_reg_7_ ( .D(wdat[7]), .C(net11820), .XR(arstz), .Q(rdat[7]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_glreg_a0_79 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module ictlr_a0 ( bkpt_ena, bkpt_pc, memaddr_c, memaddr, mcu_psr_c, mcu_psw, 
        hit_ps_c, hit_ps, mempsack, memdatao, o_set_hold, o_bkp_hold, 
        o_ofs_inc, o_inst, d_inst, sfr_psrack, sfr_psofs, sfr_psr, sfr_psw, 
        dw_rst, dw_ena, sfr_wdat, pmem_pgm, pmem_re, pmem_csb, pmem_clk, 
        pmem_a, pmem_q0, pmem_q1, pmem_twlb, wd_twlb, we_twlb, pwrdn_rst, 
        r_pwdn_en, r_multi, r_hold_mcu, clk, srst );
  input [14:0] bkpt_pc;
  input [14:0] memaddr_c;
  input [14:0] memaddr;
  input [7:0] memdatao;
  output [7:0] o_inst;
  output [7:0] d_inst;
  input [14:0] sfr_psofs;
  input [7:0] sfr_wdat;
  output [1:0] pmem_clk;
  output [15:0] pmem_a;
  input [7:0] pmem_q0;
  input [7:0] pmem_q1;
  output [1:0] pmem_twlb;
  input [1:0] wd_twlb;
  input bkpt_ena, mcu_psr_c, mcu_psw, hit_ps_c, hit_ps, sfr_psr, sfr_psw,
         dw_rst, dw_ena, we_twlb, pwrdn_rst, r_pwdn_en, r_multi, r_hold_mcu,
         clk, srst;
  output mempsack, o_set_hold, o_bkp_hold, o_ofs_inc, sfr_psrack, pmem_pgm,
         pmem_re, pmem_csb;
  wire   N152, N153, N154, N217, N218, N219, N220, N221, N222, N223, N224,
         N225, N226, N227, N228, N229, N230, N231, N232, c_buf_22__7_,
         c_buf_22__6_, c_buf_22__5_, c_buf_22__4_, c_buf_22__3_, c_buf_22__2_,
         c_buf_22__1_, c_buf_22__0_, c_buf_21__7_, c_buf_21__6_, c_buf_21__5_,
         c_buf_21__4_, c_buf_21__3_, c_buf_21__2_, c_buf_21__1_, c_buf_21__0_,
         c_buf_20__7_, c_buf_20__6_, c_buf_20__5_, c_buf_20__4_, c_buf_20__3_,
         c_buf_20__2_, c_buf_20__1_, c_buf_20__0_, c_buf_19__7_, c_buf_19__6_,
         c_buf_19__5_, c_buf_19__4_, c_buf_19__3_, c_buf_19__2_, c_buf_19__1_,
         c_buf_19__0_, c_buf_18__7_, c_buf_18__6_, c_buf_18__5_, c_buf_18__4_,
         c_buf_18__3_, c_buf_18__2_, c_buf_18__1_, c_buf_18__0_, c_buf_17__7_,
         c_buf_17__6_, c_buf_17__5_, c_buf_17__4_, c_buf_17__3_, c_buf_17__2_,
         c_buf_17__1_, c_buf_17__0_, c_buf_16__7_, c_buf_16__6_, c_buf_16__5_,
         c_buf_16__4_, c_buf_16__3_, c_buf_16__2_, c_buf_16__1_, c_buf_16__0_,
         d_psrd, r_rdy, N353, N354, N355, N356, N357, N358, N359, N431, N432,
         N433, N434, N435, N436, N437, N438, N439, N440, N441, N442, N443,
         N444, N445, N449, N450, N451, N452, N479, N480, N481, N482, N483,
         N484, N485, N486, N487, N488, N489, N490, N491, N492, N493, N494,
         N495, N496, N497, N498, N499, N500, N501, N502, N503, N504, N505,
         N506, N507, N508, N509, N510, N511, N512, N513, N514, N515, N516,
         N517, N518, N519, N520, N521, N522, N523, N524, N525, N526, N527,
         N528, N529, N530, N531, N532, N533, N534, N535, N536, N537, N538,
         N539, N540, N541, N542, N543, N544, N545, N546, N547, N548, N549,
         N550, N551, N552, N553, N554, N555, N556, N557, N558, N559, N560,
         N561, N562, N563, N564, N565, N566, N567, N568, N569, N570, N571,
         N572, N573, N574, N575, N576, N577, N578, N579, N580, N581, N582,
         N583, N584, N585, N586, N587, N588, N589, N590, N591, N592, N593,
         N594, N595, N596, N597, N598, N599, N600, N601, N602, N603, N604,
         N605, N606, N607, N608, N609, N610, N611, N612, N613, N614, N615,
         N616, N617, N618, N619, N620, N621, N622, N623, N624, N625, N626,
         N627, N628, N629, N630, N631, N632, N633, N634, N635, N636, N637,
         N638, N639, N640, N641, N642, N643, N644, N645, N646, N647, N648,
         N649, N650, N651, N652, N653, N654, N655, N656, N657, N658, N659,
         N660, N661, N662, N757, N758, N759, N786, N787, N788, N789, N790,
         N791, N792, N793, N795, N796, N797, N798, N799, N800, N801, N820,
         N821, N822, N823, N824, N825, N826, N827, N828, N829, N830, N831,
         N832, N833, N834, N835, N836, N837, N838, N839, N840, N842, N843,
         N844, N845, N846, N853, N854, N855, N856, N857, N858, N859, N860,
         N861, N862, N863, N864, N865, N866, N867, N868, N874, N875, N876,
         N877, N878, N879, N880, N881, N882, N883, N884, N885, N886, N887,
         N888, N889, N890, N891, N892, N893, N894, N895, N896, N897, N898,
         N899, cs_n, un_hold, N974, net11846, net11852, net11857, net11862,
         net11867, net11872, net11877, net11882, net11887, net11892, net11897,
         net11902, net11907, net11912, net11917, net11922, net11927, net11932,
         net11937, net11942, net11947, net11952, net11957, net11962, net11967,
         net11972, net11977, net11982, net11987, net11992, n93, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n1, n2, n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801;
  wire   [3:0] d_hold;
  wire   [1:0] dummy;
  wire   [3:0] cs_ft;
  wire   [4:0] c_ptr;
  wire   [14:0] c_adr;
  wire   [14:13] adr_p;
  wire   [7:0] rd_buf;
  wire   [7:0] dbg_01;
  wire   [7:0] dbg_02;
  wire   [7:0] dbg_03;
  wire   [7:0] dbg_04;
  wire   [7:0] dbg_05;
  wire   [7:0] dbg_06;
  wire   [7:0] dbg_07;
  wire   [7:0] dbg_08;
  wire   [7:0] dbg_09;
  wire   [7:0] dbg_0a;
  wire   [7:0] dbg_0b;
  wire   [7:0] dbg_0c;
  wire   [7:0] dbg_0d;
  wire   [7:0] dbg_0e;
  wire   [7:0] dbg_0f;
  wire   [7:0] wr_buf;
  wire   [14:0] pre_1_adr;
  wire   [6:0] wspp_cnt;
  wire   [4:0] popptr;
  wire   [4:1] sub_313_carry;
  wire   [4:2] add_255_carry;
  wire   [14:1] add_1_root_add_113_2_carry;

  DFFQX4 adr_p_reg_0_ ( .D(N854), .C(net11857), .Q(pmem_a[0]) );
  DFFQX4 adr_p_reg_1_ ( .D(N855), .C(net11857), .Q(pmem_a[1]) );
  DFFQX4 adr_p_reg_2_ ( .D(N856), .C(net11857), .Q(pmem_a[2]) );
  DFFQX4 adr_p_reg_3_ ( .D(N857), .C(net11857), .Q(pmem_a[3]) );
  DFFQX4 adr_p_reg_4_ ( .D(N858), .C(net11857), .Q(pmem_a[4]) );
  DFFQX4 adr_p_reg_5_ ( .D(N859), .C(net11857), .Q(pmem_a[5]) );
  DFFQX4 adr_p_reg_6_ ( .D(N860), .C(net11857), .Q(pmem_a[9]) );
  DFFQX4 adr_p_reg_7_ ( .D(N861), .C(net11857), .Q(pmem_a[10]) );
  DFFQX4 adr_p_reg_8_ ( .D(N862), .C(net11857), .Q(pmem_a[11]) );
  DFFQX4 adr_p_reg_9_ ( .D(N863), .C(net11857), .Q(pmem_a[12]) );
  DFFQX4 adr_p_reg_10_ ( .D(N864), .C(net11857), .Q(pmem_a[13]) );
  DFFQX4 adr_p_reg_11_ ( .D(N865), .C(net11857), .Q(pmem_a[14]) );
  DFFQX4 adr_p_reg_12_ ( .D(N866), .C(net11857), .Q(pmem_a[15]) );
  DFFQX4 a_bit_reg_0_ ( .D(N757), .C(net11852), .Q(pmem_a[6]) );
  DFFQX4 a_bit_reg_1_ ( .D(N758), .C(net11852), .Q(pmem_a[7]) );
  DFFQX4 a_bit_reg_2_ ( .D(N759), .C(net11852), .Q(pmem_a[8]) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_0 clk_gate_wspp_cnt_reg ( .CLK(clk), .EN(N899), 
        .ENCLK(net11846), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_29 clk_gate_a_bit_reg ( .CLK(clk), .EN(N898), 
        .ENCLK(net11852), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_28 clk_gate_adr_p_reg ( .CLK(clk), .EN(N853), 
        .ENCLK(net11857), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_27 clk_gate_c_buf_reg_23_ ( .CLK(clk), .EN(
        N897), .ENCLK(net11862), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_26 clk_gate_c_buf_reg_22_ ( .CLK(clk), .EN(
        N896), .ENCLK(net11867), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_25 clk_gate_c_buf_reg_21_ ( .CLK(clk), .EN(
        N895), .ENCLK(net11872), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_24 clk_gate_c_buf_reg_20_ ( .CLK(clk), .EN(
        N894), .ENCLK(net11877), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_23 clk_gate_c_buf_reg_19_ ( .CLK(clk), .EN(
        N893), .ENCLK(net11882), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_22 clk_gate_c_buf_reg_18_ ( .CLK(clk), .EN(
        N892), .ENCLK(net11887), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_21 clk_gate_c_buf_reg_17_ ( .CLK(clk), .EN(
        N891), .ENCLK(net11892), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_20 clk_gate_c_buf_reg_16_ ( .CLK(clk), .EN(
        N890), .ENCLK(net11897), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_19 clk_gate_c_buf_reg_15_ ( .CLK(clk), .EN(
        N889), .ENCLK(net11902), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_18 clk_gate_c_buf_reg_14_ ( .CLK(clk), .EN(
        N888), .ENCLK(net11907), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_17 clk_gate_c_buf_reg_13_ ( .CLK(clk), .EN(
        N887), .ENCLK(net11912), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_16 clk_gate_c_buf_reg_12_ ( .CLK(clk), .EN(
        N886), .ENCLK(net11917), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_15 clk_gate_c_buf_reg_11_ ( .CLK(clk), .EN(
        N885), .ENCLK(net11922), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_14 clk_gate_c_buf_reg_10_ ( .CLK(clk), .EN(
        N884), .ENCLK(net11927), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_13 clk_gate_c_buf_reg_9_ ( .CLK(clk), .EN(N883), .ENCLK(net11932), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_12 clk_gate_c_buf_reg_8_ ( .CLK(clk), .EN(N882), .ENCLK(net11937), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_11 clk_gate_c_buf_reg_7_ ( .CLK(clk), .EN(N881), .ENCLK(net11942), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_10 clk_gate_c_buf_reg_6_ ( .CLK(clk), .EN(N880), .ENCLK(net11947), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_9 clk_gate_c_buf_reg_5_ ( .CLK(clk), .EN(N879), 
        .ENCLK(net11952), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_8 clk_gate_c_buf_reg_4_ ( .CLK(clk), .EN(N878), 
        .ENCLK(net11957), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_7 clk_gate_c_buf_reg_3_ ( .CLK(clk), .EN(N877), 
        .ENCLK(net11962), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_6 clk_gate_c_buf_reg_2_ ( .CLK(clk), .EN(N876), 
        .ENCLK(net11967), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_5 clk_gate_c_buf_reg_1_ ( .CLK(clk), .EN(N875), 
        .ENCLK(net11972), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_4 clk_gate_c_buf_reg_0_ ( .CLK(clk), .EN(N874), 
        .ENCLK(net11977), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_3 clk_gate_c_ptr_reg ( .CLK(clk), .EN(n93), 
        .ENCLK(net11982), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_2 clk_gate_c_adr_reg ( .CLK(clk), .EN(N825), 
        .ENCLK(net11987), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_ictlr_a0_1 clk_gate_cs_ft_reg ( .CLK(clk), .EN(N820), 
        .ENCLK(net11992), .TE(1'b0) );
  ictlr_a0_DW01_inc_1 add_242 ( .A(c_adr), .SUM({N445, N444, N443, N442, N441, 
        N440, N439, N438, N437, N436, N435, N434, N433, N432, N431}) );
  ictlr_a0_DW01_inc_2 r492 ( .A({adr_p, pmem_a[15:9], pmem_a[5:0]}), .SUM(
        pre_1_adr) );
  FAD1X1 sub_313_U2_1 ( .A(memaddr[1]), .B(n430), .CI(sub_313_carry[1]), .CO(
        sub_313_carry[2]), .SO(popptr[1]) );
  FAD1X1 sub_313_U2_2 ( .A(memaddr[2]), .B(n119), .CI(sub_313_carry[2]), .CO(
        sub_313_carry[3]), .SO(popptr[2]) );
  FAD1X1 sub_313_U2_3 ( .A(memaddr[3]), .B(n431), .CI(sub_313_carry[3]), .CO(
        sub_313_carry[4]), .SO(popptr[3]) );
  HAD1X1 add_255_U1_1_1 ( .A(c_ptr[1]), .B(c_ptr[0]), .CO(add_255_carry[2]), 
        .SO(N449) );
  HAD1X1 add_255_U1_1_2 ( .A(c_ptr[2]), .B(add_255_carry[2]), .CO(
        add_255_carry[3]), .SO(N450) );
  HAD1X1 add_255_U1_1_3 ( .A(c_ptr[3]), .B(add_255_carry[3]), .CO(
        add_255_carry[4]), .SO(N451) );
  FAD1X1 add_1_root_add_113_2_U1_1 ( .A(c_adr[1]), .B(c_ptr[1]), .CI(
        add_1_root_add_113_2_carry[1]), .CO(add_1_root_add_113_2_carry[2]), 
        .SO(N218) );
  FAD1X1 add_1_root_add_113_2_U1_2 ( .A(c_adr[2]), .B(c_ptr[2]), .CI(
        add_1_root_add_113_2_carry[2]), .CO(add_1_root_add_113_2_carry[3]), 
        .SO(N219) );
  FAD1X1 add_1_root_add_113_2_U1_3 ( .A(c_adr[3]), .B(c_ptr[3]), .CI(
        add_1_root_add_113_2_carry[3]), .CO(add_1_root_add_113_2_carry[4]), 
        .SO(N220) );
  FAD1X1 add_1_root_add_113_2_U1_4 ( .A(c_adr[4]), .B(c_ptr[4]), .CI(
        add_1_root_add_113_2_carry[4]), .CO(add_1_root_add_113_2_carry[5]), 
        .SO(N221) );
  DFFQX1 wspp_cnt_reg_1_ ( .D(N796), .C(net11846), .Q(wspp_cnt[1]) );
  DFFQX1 wspp_cnt_reg_2_ ( .D(N797), .C(net11846), .Q(wspp_cnt[2]) );
  DFFQX1 wspp_cnt_reg_0_ ( .D(N795), .C(net11846), .Q(wspp_cnt[0]) );
  DFFQX1 d_hold_reg_3_ ( .D(N154), .C(clk), .Q(d_hold[3]) );
  DFFQX1 dummy_reg_1_ ( .D(n650), .C(clk), .Q(dummy[1]) );
  DFFQX1 d_hold_reg_1_ ( .D(N152), .C(clk), .Q(d_hold[1]) );
  DFFQX1 d_hold_reg_2_ ( .D(N153), .C(clk), .Q(d_hold[2]) );
  DFFQX1 dummy_reg_0_ ( .D(n651), .C(clk), .Q(dummy[0]) );
  DFFQX1 d_hold_reg_0_ ( .D(n801), .C(clk), .Q(d_hold[0]) );
  DFFQX1 d_psrd_reg ( .D(n649), .C(net11992), .Q(d_psrd) );
  DFFQX1 c_adr_reg_14_ ( .D(N840), .C(net11987), .Q(c_adr[14]) );
  DFFQX1 c_adr_reg_12_ ( .D(N838), .C(net11987), .Q(c_adr[12]) );
  DFFQX1 c_adr_reg_13_ ( .D(N839), .C(net11987), .Q(c_adr[13]) );
  DFFQX1 c_adr_reg_11_ ( .D(N837), .C(net11987), .Q(c_adr[11]) );
  DFFQX1 c_adr_reg_8_ ( .D(N834), .C(net11987), .Q(c_adr[8]) );
  DFFQX1 c_adr_reg_9_ ( .D(N835), .C(net11987), .Q(c_adr[9]) );
  DFFQX1 c_adr_reg_10_ ( .D(N836), .C(net11987), .Q(c_adr[10]) );
  DFFQX1 c_adr_reg_6_ ( .D(N832), .C(net11987), .Q(c_adr[6]) );
  DFFQX1 c_adr_reg_7_ ( .D(N833), .C(net11987), .Q(c_adr[7]) );
  DFFQX1 c_adr_reg_5_ ( .D(N831), .C(net11987), .Q(c_adr[5]) );
  DFFQX1 c_ptr_reg_4_ ( .D(N846), .C(net11982), .Q(c_ptr[4]) );
  DFFQX1 c_ptr_reg_2_ ( .D(N844), .C(net11982), .Q(c_ptr[2]) );
  DFFQX1 c_ptr_reg_3_ ( .D(N845), .C(net11982), .Q(c_ptr[3]) );
  DFFQX1 c_ptr_reg_0_ ( .D(N842), .C(net11982), .Q(c_ptr[0]) );
  DFFQX1 c_ptr_reg_1_ ( .D(N843), .C(net11982), .Q(c_ptr[1]) );
  DFFQX1 pgm_p_reg ( .D(n644), .C(net11992), .Q(pmem_pgm) );
  DFFQX1 un_hold_reg ( .D(N974), .C(clk), .Q(un_hold) );
  DFFQX1 c_buf_reg_5__6_ ( .D(N525), .C(net11952), .Q(dbg_05[6]) );
  DFFQX1 c_buf_reg_2__6_ ( .D(N501), .C(net11967), .Q(dbg_02[6]) );
  DFFQX1 c_buf_reg_5__4_ ( .D(N523), .C(net11952), .Q(dbg_05[4]) );
  DFFQX1 c_buf_reg_2__4_ ( .D(N499), .C(net11967), .Q(dbg_02[4]) );
  DFFQX1 c_buf_reg_5__3_ ( .D(N522), .C(net11952), .Q(dbg_05[3]) );
  DFFQX1 c_buf_reg_2__3_ ( .D(N498), .C(net11967), .Q(dbg_02[3]) );
  DFFQX1 c_buf_reg_5__2_ ( .D(N521), .C(net11952), .Q(dbg_05[2]) );
  DFFQX1 c_buf_reg_2__2_ ( .D(N497), .C(net11967), .Q(dbg_02[2]) );
  DFFQX1 c_buf_reg_5__1_ ( .D(N520), .C(net11952), .Q(dbg_05[1]) );
  DFFQX1 c_buf_reg_2__1_ ( .D(N496), .C(net11967), .Q(dbg_02[1]) );
  DFFQX1 c_buf_reg_5__0_ ( .D(N519), .C(net11952), .Q(dbg_05[0]) );
  DFFQX1 c_buf_reg_2__0_ ( .D(N495), .C(net11967), .Q(dbg_02[0]) );
  DFFQX1 c_buf_reg_3__6_ ( .D(N509), .C(net11962), .Q(dbg_03[6]) );
  DFFQX1 c_buf_reg_3__5_ ( .D(N508), .C(net11962), .Q(dbg_03[5]) );
  DFFQX1 c_buf_reg_3__4_ ( .D(N507), .C(net11962), .Q(dbg_03[4]) );
  DFFQX1 c_buf_reg_3__3_ ( .D(N506), .C(net11962), .Q(dbg_03[3]) );
  DFFQX1 c_buf_reg_3__2_ ( .D(N505), .C(net11962), .Q(dbg_03[2]) );
  DFFQX1 c_buf_reg_3__1_ ( .D(N504), .C(net11962), .Q(dbg_03[1]) );
  DFFQX1 c_buf_reg_3__0_ ( .D(N503), .C(net11962), .Q(dbg_03[0]) );
  DFFQX1 c_buf_reg_4__6_ ( .D(N517), .C(net11957), .Q(dbg_04[6]) );
  DFFQX1 c_buf_reg_1__6_ ( .D(N493), .C(net11972), .Q(dbg_01[6]) );
  DFFQX1 c_buf_reg_4__4_ ( .D(N515), .C(net11957), .Q(dbg_04[4]) );
  DFFQX1 c_buf_reg_1__4_ ( .D(N491), .C(net11972), .Q(dbg_01[4]) );
  DFFQX1 c_buf_reg_4__3_ ( .D(N514), .C(net11957), .Q(dbg_04[3]) );
  DFFQX1 c_buf_reg_1__3_ ( .D(N490), .C(net11972), .Q(dbg_01[3]) );
  DFFQX1 c_buf_reg_4__2_ ( .D(N513), .C(net11957), .Q(dbg_04[2]) );
  DFFQX1 c_buf_reg_1__2_ ( .D(N489), .C(net11972), .Q(dbg_01[2]) );
  DFFQX1 c_buf_reg_4__1_ ( .D(N512), .C(net11957), .Q(dbg_04[1]) );
  DFFQX1 c_buf_reg_1__1_ ( .D(N488), .C(net11972), .Q(dbg_01[1]) );
  DFFQX1 c_buf_reg_4__0_ ( .D(N511), .C(net11957), .Q(dbg_04[0]) );
  DFFQX1 c_buf_reg_1__0_ ( .D(N487), .C(net11972), .Q(dbg_01[0]) );
  DFFQX1 c_buf_reg_0__6_ ( .D(N485), .C(net11977), .Q(rd_buf[6]) );
  DFFQX1 c_buf_reg_0__5_ ( .D(N484), .C(net11977), .Q(rd_buf[5]) );
  DFFQX1 c_buf_reg_0__3_ ( .D(N482), .C(net11977), .Q(rd_buf[3]) );
  DFFQX1 c_buf_reg_0__2_ ( .D(N481), .C(net11977), .Q(rd_buf[2]) );
  DFFQX1 c_buf_reg_0__1_ ( .D(N480), .C(net11977), .Q(rd_buf[1]) );
  DFFQX1 c_buf_reg_6__6_ ( .D(N533), .C(net11947), .Q(dbg_06[6]) );
  DFFQX1 c_buf_reg_6__5_ ( .D(N532), .C(net11947), .Q(dbg_06[5]) );
  DFFQX1 c_buf_reg_6__4_ ( .D(N531), .C(net11947), .Q(dbg_06[4]) );
  DFFQX1 c_buf_reg_6__3_ ( .D(N530), .C(net11947), .Q(dbg_06[3]) );
  DFFQX1 c_buf_reg_6__2_ ( .D(N529), .C(net11947), .Q(dbg_06[2]) );
  DFFQX1 c_buf_reg_6__1_ ( .D(N528), .C(net11947), .Q(dbg_06[1]) );
  DFFQX1 c_buf_reg_6__0_ ( .D(N527), .C(net11947), .Q(dbg_06[0]) );
  DFFQX1 c_buf_reg_0__4_ ( .D(N483), .C(net11977), .Q(rd_buf[4]) );
  DFFQX1 c_buf_reg_0__0_ ( .D(N479), .C(net11977), .Q(rd_buf[0]) );
  DFFQX1 re_p_reg ( .D(n647), .C(clk), .Q(pmem_re) );
  DFFQX1 c_buf_reg_11__4_ ( .D(N571), .C(net11922), .Q(dbg_0b[4]) );
  DFFQX1 c_buf_reg_11__3_ ( .D(N570), .C(net11922), .Q(dbg_0b[3]) );
  DFFQX1 c_buf_reg_11__2_ ( .D(N569), .C(net11922), .Q(dbg_0b[2]) );
  DFFQX1 c_buf_reg_11__1_ ( .D(N568), .C(net11922), .Q(dbg_0b[1]) );
  DFFQX1 c_buf_reg_11__0_ ( .D(N567), .C(net11922), .Q(dbg_0b[0]) );
  DFFQX1 c_buf_reg_10__6_ ( .D(N565), .C(net11927), .Q(dbg_0a[6]) );
  DFFQX1 c_buf_reg_10__4_ ( .D(N563), .C(net11927), .Q(dbg_0a[4]) );
  DFFQX1 c_buf_reg_10__3_ ( .D(N562), .C(net11927), .Q(dbg_0a[3]) );
  DFFQX1 c_buf_reg_10__2_ ( .D(N561), .C(net11927), .Q(dbg_0a[2]) );
  DFFQX1 c_buf_reg_10__1_ ( .D(N560), .C(net11927), .Q(dbg_0a[1]) );
  DFFQX1 c_buf_reg_10__0_ ( .D(N559), .C(net11927), .Q(dbg_0a[0]) );
  DFFQX1 c_buf_reg_7__4_ ( .D(N539), .C(net11942), .Q(dbg_07[4]) );
  DFFQX1 c_buf_reg_5__5_ ( .D(N524), .C(net11952), .Q(dbg_05[5]) );
  DFFQX1 c_buf_reg_2__5_ ( .D(N500), .C(net11967), .Q(dbg_02[5]) );
  DFFQX1 c_buf_reg_4__5_ ( .D(N516), .C(net11957), .Q(dbg_04[5]) );
  DFFQX1 c_buf_reg_1__5_ ( .D(N492), .C(net11972), .Q(dbg_01[5]) );
  DFFQX1 r_twlb_reg_0_ ( .D(n646), .C(clk), .Q(pmem_twlb[0]) );
  DFFQX1 adr_p_reg_14_ ( .D(N868), .C(net11857), .Q(adr_p[14]) );
  DFFQX1 c_buf_reg_22__6_ ( .D(N661), .C(net11867), .Q(c_buf_22__6_) );
  DFFQX1 c_buf_reg_22__4_ ( .D(N659), .C(net11867), .Q(c_buf_22__4_) );
  DFFQX1 c_buf_reg_22__3_ ( .D(N658), .C(net11867), .Q(c_buf_22__3_) );
  DFFQX1 c_buf_reg_22__2_ ( .D(N657), .C(net11867), .Q(c_buf_22__2_) );
  DFFQX1 c_buf_reg_22__1_ ( .D(N656), .C(net11867), .Q(c_buf_22__1_) );
  DFFQX1 c_buf_reg_22__0_ ( .D(N655), .C(net11867), .Q(c_buf_22__0_) );
  DFFQX1 c_buf_reg_21__6_ ( .D(N653), .C(net11872), .Q(c_buf_21__6_) );
  DFFQX1 c_buf_reg_21__4_ ( .D(N651), .C(net11872), .Q(c_buf_21__4_) );
  DFFQX1 c_buf_reg_21__3_ ( .D(N650), .C(net11872), .Q(c_buf_21__3_) );
  DFFQX1 c_buf_reg_21__2_ ( .D(N649), .C(net11872), .Q(c_buf_21__2_) );
  DFFQX1 c_buf_reg_21__1_ ( .D(N648), .C(net11872), .Q(c_buf_21__1_) );
  DFFQX1 c_buf_reg_21__0_ ( .D(N647), .C(net11872), .Q(c_buf_21__0_) );
  DFFQX1 c_buf_reg_20__6_ ( .D(N645), .C(net11877), .Q(c_buf_20__6_) );
  DFFQX1 c_buf_reg_20__5_ ( .D(N644), .C(net11877), .Q(c_buf_20__5_) );
  DFFQX1 c_buf_reg_20__4_ ( .D(N643), .C(net11877), .Q(c_buf_20__4_) );
  DFFQX1 c_buf_reg_20__3_ ( .D(N642), .C(net11877), .Q(c_buf_20__3_) );
  DFFQX1 c_buf_reg_20__2_ ( .D(N641), .C(net11877), .Q(c_buf_20__2_) );
  DFFQX1 c_buf_reg_20__1_ ( .D(N640), .C(net11877), .Q(c_buf_20__1_) );
  DFFQX1 c_buf_reg_20__0_ ( .D(N639), .C(net11877), .Q(c_buf_20__0_) );
  DFFQX1 c_buf_reg_19__6_ ( .D(N637), .C(net11882), .Q(c_buf_19__6_) );
  DFFQX1 c_buf_reg_19__4_ ( .D(N635), .C(net11882), .Q(c_buf_19__4_) );
  DFFQX1 c_buf_reg_19__3_ ( .D(N634), .C(net11882), .Q(c_buf_19__3_) );
  DFFQX1 c_buf_reg_19__2_ ( .D(N633), .C(net11882), .Q(c_buf_19__2_) );
  DFFQX1 c_buf_reg_19__1_ ( .D(N632), .C(net11882), .Q(c_buf_19__1_) );
  DFFQX1 c_buf_reg_19__0_ ( .D(N631), .C(net11882), .Q(c_buf_19__0_) );
  DFFQX1 c_buf_reg_18__6_ ( .D(N629), .C(net11887), .Q(c_buf_18__6_) );
  DFFQX1 c_buf_reg_18__4_ ( .D(N627), .C(net11887), .Q(c_buf_18__4_) );
  DFFQX1 c_buf_reg_18__3_ ( .D(N626), .C(net11887), .Q(c_buf_18__3_) );
  DFFQX1 c_buf_reg_18__2_ ( .D(N625), .C(net11887), .Q(c_buf_18__2_) );
  DFFQX1 c_buf_reg_18__1_ ( .D(N624), .C(net11887), .Q(c_buf_18__1_) );
  DFFQX1 c_buf_reg_18__0_ ( .D(N623), .C(net11887), .Q(c_buf_18__0_) );
  DFFQX1 c_buf_reg_17__6_ ( .D(N621), .C(net11892), .Q(c_buf_17__6_) );
  DFFQX1 c_buf_reg_17__5_ ( .D(N620), .C(net11892), .Q(c_buf_17__5_) );
  DFFQX1 c_buf_reg_17__4_ ( .D(N619), .C(net11892), .Q(c_buf_17__4_) );
  DFFQX1 c_buf_reg_17__3_ ( .D(N618), .C(net11892), .Q(c_buf_17__3_) );
  DFFQX1 c_buf_reg_17__2_ ( .D(N617), .C(net11892), .Q(c_buf_17__2_) );
  DFFQX1 c_buf_reg_17__1_ ( .D(N616), .C(net11892), .Q(c_buf_17__1_) );
  DFFQX1 c_buf_reg_17__0_ ( .D(N615), .C(net11892), .Q(c_buf_17__0_) );
  DFFQX1 c_buf_reg_16__6_ ( .D(N613), .C(net11897), .Q(c_buf_16__6_) );
  DFFQX1 c_buf_reg_16__4_ ( .D(N611), .C(net11897), .Q(c_buf_16__4_) );
  DFFQX1 c_buf_reg_16__3_ ( .D(N610), .C(net11897), .Q(c_buf_16__3_) );
  DFFQX1 c_buf_reg_16__2_ ( .D(N609), .C(net11897), .Q(c_buf_16__2_) );
  DFFQX1 c_buf_reg_16__1_ ( .D(N608), .C(net11897), .Q(c_buf_16__1_) );
  DFFQX1 c_buf_reg_16__0_ ( .D(N607), .C(net11897), .Q(c_buf_16__0_) );
  DFFQX1 c_buf_reg_15__6_ ( .D(N605), .C(net11902), .Q(dbg_0f[6]) );
  DFFQX1 c_buf_reg_15__5_ ( .D(N604), .C(net11902), .Q(dbg_0f[5]) );
  DFFQX1 c_buf_reg_15__4_ ( .D(N603), .C(net11902), .Q(dbg_0f[4]) );
  DFFQX1 c_buf_reg_15__3_ ( .D(N602), .C(net11902), .Q(dbg_0f[3]) );
  DFFQX1 c_buf_reg_15__2_ ( .D(N601), .C(net11902), .Q(dbg_0f[2]) );
  DFFQX1 c_buf_reg_15__1_ ( .D(N600), .C(net11902), .Q(dbg_0f[1]) );
  DFFQX1 c_buf_reg_15__0_ ( .D(N599), .C(net11902), .Q(dbg_0f[0]) );
  DFFQX1 c_buf_reg_14__6_ ( .D(N597), .C(net11907), .Q(dbg_0e[6]) );
  DFFQX1 c_buf_reg_14__5_ ( .D(N596), .C(net11907), .Q(dbg_0e[5]) );
  DFFQX1 c_buf_reg_14__4_ ( .D(N595), .C(net11907), .Q(dbg_0e[4]) );
  DFFQX1 c_buf_reg_14__3_ ( .D(N594), .C(net11907), .Q(dbg_0e[3]) );
  DFFQX1 c_buf_reg_14__2_ ( .D(N593), .C(net11907), .Q(dbg_0e[2]) );
  DFFQX1 c_buf_reg_14__1_ ( .D(N592), .C(net11907), .Q(dbg_0e[1]) );
  DFFQX1 c_buf_reg_14__0_ ( .D(N591), .C(net11907), .Q(dbg_0e[0]) );
  DFFQX1 c_buf_reg_13__6_ ( .D(N589), .C(net11912), .Q(dbg_0d[6]) );
  DFFQX1 c_buf_reg_13__5_ ( .D(N588), .C(net11912), .Q(dbg_0d[5]) );
  DFFQX1 c_buf_reg_13__4_ ( .D(N587), .C(net11912), .Q(dbg_0d[4]) );
  DFFQX1 c_buf_reg_13__3_ ( .D(N586), .C(net11912), .Q(dbg_0d[3]) );
  DFFQX1 c_buf_reg_13__2_ ( .D(N585), .C(net11912), .Q(dbg_0d[2]) );
  DFFQX1 c_buf_reg_13__1_ ( .D(N584), .C(net11912), .Q(dbg_0d[1]) );
  DFFQX1 c_buf_reg_13__0_ ( .D(N583), .C(net11912), .Q(dbg_0d[0]) );
  DFFQX1 c_buf_reg_12__6_ ( .D(N581), .C(net11917), .Q(dbg_0c[6]) );
  DFFQX1 c_buf_reg_12__5_ ( .D(N580), .C(net11917), .Q(dbg_0c[5]) );
  DFFQX1 c_buf_reg_12__4_ ( .D(N579), .C(net11917), .Q(dbg_0c[4]) );
  DFFQX1 c_buf_reg_12__3_ ( .D(N578), .C(net11917), .Q(dbg_0c[3]) );
  DFFQX1 c_buf_reg_12__2_ ( .D(N577), .C(net11917), .Q(dbg_0c[2]) );
  DFFQX1 c_buf_reg_12__1_ ( .D(N576), .C(net11917), .Q(dbg_0c[1]) );
  DFFQX1 c_buf_reg_12__0_ ( .D(N575), .C(net11917), .Q(dbg_0c[0]) );
  DFFQX1 c_buf_reg_11__6_ ( .D(N573), .C(net11922), .Q(dbg_0b[6]) );
  DFFQX1 c_buf_reg_11__5_ ( .D(N572), .C(net11922), .Q(dbg_0b[5]) );
  DFFQX1 c_buf_reg_10__5_ ( .D(N564), .C(net11927), .Q(dbg_0a[5]) );
  DFFQX1 c_buf_reg_9__6_ ( .D(N557), .C(net11932), .Q(dbg_09[6]) );
  DFFQX1 c_buf_reg_9__5_ ( .D(N556), .C(net11932), .Q(dbg_09[5]) );
  DFFQX1 c_buf_reg_9__4_ ( .D(N555), .C(net11932), .Q(dbg_09[4]) );
  DFFQX1 c_buf_reg_9__3_ ( .D(N554), .C(net11932), .Q(dbg_09[3]) );
  DFFQX1 c_buf_reg_9__2_ ( .D(N553), .C(net11932), .Q(dbg_09[2]) );
  DFFQX1 c_buf_reg_9__1_ ( .D(N552), .C(net11932), .Q(dbg_09[1]) );
  DFFQX1 c_buf_reg_9__0_ ( .D(N551), .C(net11932), .Q(dbg_09[0]) );
  DFFQX1 c_buf_reg_8__6_ ( .D(N549), .C(net11937), .Q(dbg_08[6]) );
  DFFQX1 c_buf_reg_8__5_ ( .D(N548), .C(net11937), .Q(dbg_08[5]) );
  DFFQX1 c_buf_reg_8__4_ ( .D(N547), .C(net11937), .Q(dbg_08[4]) );
  DFFQX1 c_buf_reg_8__3_ ( .D(N546), .C(net11937), .Q(dbg_08[3]) );
  DFFQX1 c_buf_reg_8__2_ ( .D(N545), .C(net11937), .Q(dbg_08[2]) );
  DFFQX1 c_buf_reg_8__1_ ( .D(N544), .C(net11937), .Q(dbg_08[1]) );
  DFFQX1 c_buf_reg_8__0_ ( .D(N543), .C(net11937), .Q(dbg_08[0]) );
  DFFQX1 c_buf_reg_7__6_ ( .D(N541), .C(net11942), .Q(dbg_07[6]) );
  DFFQX1 c_buf_reg_7__5_ ( .D(N540), .C(net11942), .Q(dbg_07[5]) );
  DFFQX1 c_buf_reg_7__3_ ( .D(N538), .C(net11942), .Q(dbg_07[3]) );
  DFFQX1 c_buf_reg_7__2_ ( .D(N537), .C(net11942), .Q(dbg_07[2]) );
  DFFQX1 c_buf_reg_7__1_ ( .D(N536), .C(net11942), .Q(dbg_07[1]) );
  DFFQX1 c_buf_reg_7__0_ ( .D(N535), .C(net11942), .Q(dbg_07[0]) );
  DFFQX1 c_buf_reg_23__4_ ( .D(N790), .C(net11862), .Q(wr_buf[4]) );
  DFFQX1 c_buf_reg_23__6_ ( .D(N792), .C(net11862), .Q(wr_buf[6]) );
  DFFQX1 c_buf_reg_23__2_ ( .D(N788), .C(net11862), .Q(wr_buf[2]) );
  DFFQX1 c_buf_reg_23__3_ ( .D(N789), .C(net11862), .Q(wr_buf[3]) );
  DFFQX1 c_buf_reg_23__5_ ( .D(N791), .C(net11862), .Q(wr_buf[5]) );
  DFFQX1 c_buf_reg_23__1_ ( .D(N787), .C(net11862), .Q(wr_buf[1]) );
  DFFQX1 c_buf_reg_23__0_ ( .D(N786), .C(net11862), .Q(wr_buf[0]) );
  DFFQX1 adr_p_reg_13_ ( .D(N867), .C(net11857), .Q(adr_p[13]) );
  DFFQX1 c_buf_reg_5__7_ ( .D(N526), .C(net11952), .Q(dbg_05[7]) );
  DFFQX1 c_buf_reg_2__7_ ( .D(N502), .C(net11967), .Q(dbg_02[7]) );
  DFFQX1 c_buf_reg_3__7_ ( .D(N510), .C(net11962), .Q(dbg_03[7]) );
  DFFQX1 c_buf_reg_4__7_ ( .D(N518), .C(net11957), .Q(dbg_04[7]) );
  DFFQX1 c_buf_reg_1__7_ ( .D(N494), .C(net11972), .Q(dbg_01[7]) );
  DFFQX1 c_buf_reg_0__7_ ( .D(N486), .C(net11977), .Q(rd_buf[7]) );
  DFFQX1 c_buf_reg_6__7_ ( .D(N534), .C(net11947), .Q(dbg_06[7]) );
  DFFQX1 r_twlb_reg_1_ ( .D(n645), .C(clk), .Q(pmem_twlb[1]) );
  DFFQX1 wspp_cnt_reg_5_ ( .D(N800), .C(net11846), .Q(wspp_cnt[5]) );
  DFFQX1 wspp_cnt_reg_3_ ( .D(N798), .C(net11846), .Q(wspp_cnt[3]) );
  DFFQX1 wspp_cnt_reg_4_ ( .D(N799), .C(net11846), .Q(wspp_cnt[4]) );
  DFFQX1 wspp_cnt_reg_6_ ( .D(N801), .C(net11846), .Q(wspp_cnt[6]) );
  DFFQX1 c_buf_reg_22__5_ ( .D(N660), .C(net11867), .Q(c_buf_22__5_) );
  DFFQX1 c_buf_reg_21__5_ ( .D(N652), .C(net11872), .Q(c_buf_21__5_) );
  DFFQX1 c_buf_reg_19__5_ ( .D(N636), .C(net11882), .Q(c_buf_19__5_) );
  DFFQX1 c_buf_reg_18__5_ ( .D(N628), .C(net11887), .Q(c_buf_18__5_) );
  DFFQX1 c_buf_reg_16__5_ ( .D(N612), .C(net11897), .Q(c_buf_16__5_) );
  DFFQX1 c_buf_reg_14__7_ ( .D(N598), .C(net11907), .Q(dbg_0e[7]) );
  DFFQX1 c_buf_reg_11__7_ ( .D(N574), .C(net11922), .Q(dbg_0b[7]) );
  DFFQX1 c_buf_reg_10__7_ ( .D(N566), .C(net11927), .Q(dbg_0a[7]) );
  DFFQX1 c_buf_reg_8__7_ ( .D(N550), .C(net11937), .Q(dbg_08[7]) );
  DFFQX1 c_buf_reg_7__7_ ( .D(N542), .C(net11942), .Q(dbg_07[7]) );
  DFFQX1 c_buf_reg_22__7_ ( .D(N662), .C(net11867), .Q(c_buf_22__7_) );
  DFFQX1 c_buf_reg_21__7_ ( .D(N654), .C(net11872), .Q(c_buf_21__7_) );
  DFFQX1 c_buf_reg_20__7_ ( .D(N646), .C(net11877), .Q(c_buf_20__7_) );
  DFFQX1 c_buf_reg_19__7_ ( .D(N638), .C(net11882), .Q(c_buf_19__7_) );
  DFFQX1 c_buf_reg_18__7_ ( .D(N630), .C(net11887), .Q(c_buf_18__7_) );
  DFFQX1 c_buf_reg_17__7_ ( .D(N622), .C(net11892), .Q(c_buf_17__7_) );
  DFFQX1 c_buf_reg_16__7_ ( .D(N614), .C(net11897), .Q(c_buf_16__7_) );
  DFFQX1 c_buf_reg_15__7_ ( .D(N606), .C(net11902), .Q(dbg_0f[7]) );
  DFFQX1 c_buf_reg_13__7_ ( .D(N590), .C(net11912), .Q(dbg_0d[7]) );
  DFFQX1 c_buf_reg_12__7_ ( .D(N582), .C(net11917), .Q(dbg_0c[7]) );
  DFFQX1 c_buf_reg_9__7_ ( .D(N558), .C(net11932), .Q(dbg_09[7]) );
  DFFQX1 c_buf_reg_23__7_ ( .D(N793), .C(net11862), .Q(wr_buf[7]) );
  DFFQX1 r_rdy_reg ( .D(n648), .C(clk), .Q(r_rdy) );
  DFFQX1 cs_ft_reg_2_ ( .D(N823), .C(net11992), .Q(cs_ft[2]) );
  DFFQX1 cs_ft_reg_3_ ( .D(N824), .C(net11992), .Q(cs_ft[3]) );
  DFFQX1 cs_ft_reg_1_ ( .D(N822), .C(net11992), .Q(cs_ft[1]) );
  DFFQX1 cs_ft_reg_0_ ( .D(N821), .C(net11992), .Q(cs_ft[0]) );
  DFFQX1 c_adr_reg_3_ ( .D(N829), .C(net11987), .Q(c_adr[3]) );
  DFFQX1 c_adr_reg_4_ ( .D(N830), .C(net11987), .Q(c_adr[4]) );
  DFFQX1 c_adr_reg_2_ ( .D(N828), .C(net11987), .Q(c_adr[2]) );
  DFFQX1 c_adr_reg_0_ ( .D(N826), .C(net11987), .Q(c_adr[0]) );
  DFFQX1 c_adr_reg_1_ ( .D(N827), .C(net11987), .Q(c_adr[1]) );
  DFFNQXL ck_n_reg_0_ ( .D(n641), .XC(clk), .Q(pmem_clk[0]) );
  DFFNQXL cs_n_reg ( .D(n643), .XC(clk), .Q(cs_n) );
  DFFNQXL ck_n_reg_1_ ( .D(n642), .XC(clk), .Q(pmem_clk[1]) );
  XOR3X1 sub_313_U2_4 ( .A(memaddr[4]), .B(n432), .C(sub_313_carry[4]), .Y(
        popptr[4]) );
  INVX1 U3 ( .A(n120), .Y(n121) );
  OA222X1 U4 ( .A(memaddr_c[4]), .B(n62), .C(n165), .D(n164), .E(memaddr_c[5]), 
        .F(n64), .Y(n170) );
  OAI211X1 U5 ( .C(n437), .D(n122), .A(n121), .B(n436), .Y(n123) );
  NOR3XL U6 ( .A(n367), .B(n65), .C(n273), .Y(n40) );
  NAND21X1 U7 ( .B(n199), .A(n198), .Y(n374) );
  OA22X1 U8 ( .A(n399), .B(n2), .C(n400), .D(n196), .Y(n1) );
  INVX1 U9 ( .A(n379), .Y(n301) );
  XNOR2XL U10 ( .A(n147), .B(c_adr[14]), .Y(n2) );
  INVXL U11 ( .A(n343), .Y(n3) );
  INVXL U12 ( .A(n3), .Y(n4) );
  INVX1 U13 ( .A(n292), .Y(n5) );
  INVX1 U14 ( .A(n292), .Y(n6) );
  INVX1 U15 ( .A(n290), .Y(n7) );
  INVX1 U16 ( .A(n290), .Y(n8) );
  INVX1 U17 ( .A(n289), .Y(n9) );
  INVX1 U18 ( .A(n289), .Y(n10) );
  INVX1 U19 ( .A(n288), .Y(n11) );
  INVX1 U20 ( .A(n288), .Y(n12) );
  INVX1 U21 ( .A(n287), .Y(n13) );
  INVX1 U22 ( .A(n287), .Y(n14) );
  INVX1 U23 ( .A(n340), .Y(n15) );
  BUFX3 U24 ( .A(n358), .Y(n16) );
  INVX1 U25 ( .A(n286), .Y(n17) );
  INVX1 U26 ( .A(n286), .Y(n18) );
  INVX1 U27 ( .A(n736), .Y(n19) );
  INVX1 U28 ( .A(n266), .Y(n20) );
  INVX1 U29 ( .A(n320), .Y(n21) );
  INVX1 U30 ( .A(n285), .Y(n22) );
  INVX1 U31 ( .A(n285), .Y(n23) );
  INVX1 U32 ( .A(n318), .Y(n24) );
  INVX1 U33 ( .A(n415), .Y(n25) );
  NAND21X1 U34 ( .B(d_psrd), .A(n232), .Y(n379) );
  INVXL U35 ( .A(n87), .Y(n26) );
  INVXL U36 ( .A(n87), .Y(n27) );
  OAI32X1 U37 ( .A(n389), .B(d_psrd), .C(n85), .D(n376), .E(n312), .Y(n344) );
  INVXL U38 ( .A(n315), .Y(n28) );
  INVXL U39 ( .A(n315), .Y(n29) );
  INVX1 U40 ( .A(n284), .Y(n30) );
  INVX1 U41 ( .A(n284), .Y(n31) );
  NAND21X1 U42 ( .B(pwrdn_rst), .A(n88), .Y(n382) );
  GEN2XL U43 ( .D(n280), .E(n279), .C(n278), .B(n86), .A(n277), .Y(n642) );
  INVX1 U44 ( .A(n379), .Y(n66) );
  OAI222XL U45 ( .A(memaddr_c[13]), .B(n195), .C(n194), .D(n193), .E(
        memaddr_c[12]), .F(n192), .Y(n33) );
  GEN2XL U46 ( .D(n280), .E(n275), .C(n278), .B(n87), .A(n274), .Y(n641) );
  INVX1 U47 ( .A(n349), .Y(n232) );
  NAND2X1 U48 ( .A(n343), .B(pre_1_adr[14]), .Y(n333) );
  INVXL U49 ( .A(n315), .Y(n260) );
  NAND2XL U50 ( .A(n87), .B(n395), .Y(n322) );
  AND2XL U51 ( .A(n87), .B(n316), .Y(n37) );
  OA21XL U52 ( .B(n413), .C(n211), .A(n210), .Y(n226) );
  NAND21XL U53 ( .B(n726), .A(n66), .Y(n266) );
  INVXL U54 ( .A(memaddr_c[1]), .Y(n412) );
  NAND31XL U55 ( .C(n325), .A(n32), .B(n315), .Y(N897) );
  AOI21X1 U56 ( .B(n265), .C(n264), .A(n263), .Y(n32) );
  INVXL U57 ( .A(n227), .Y(n160) );
  INVXL U58 ( .A(n301), .Y(n84) );
  INVXL U59 ( .A(memaddr_c[0]), .Y(n413) );
  OAI32XL U60 ( .A(n171), .B(n170), .C(n169), .D(memaddr_c[6]), .E(n168), .Y(
        n172) );
  AO21XL U61 ( .B(memaddr_c[6]), .C(n143), .A(n117), .Y(n120) );
  OAI21BBX1 U62 ( .A(n183), .B(n182), .C(n220), .Y(n185) );
  AOI21XL U63 ( .B(n16), .C(memaddr_c[6]), .A(n26), .Y(n44) );
  NAND2X1 U64 ( .A(n33), .B(n1), .Y(n213) );
  NAND32X1 U65 ( .B(n276), .C(n240), .A(n229), .Y(n303) );
  OAI21BBX1 U66 ( .A(n163), .B(n162), .C(n218), .Y(n164) );
  INVX1 U67 ( .A(n374), .Y(n233) );
  INVXL U68 ( .A(memaddr_c[6]), .Y(n407) );
  AND3X1 U69 ( .A(pmem_clk[1]), .B(n40), .C(n276), .Y(n277) );
  AOI21XL U70 ( .B(n16), .C(memaddr_c[0]), .A(n27), .Y(n58) );
  OAI21BBX1 U71 ( .A(n339), .B(n338), .C(n34), .Y(n645) );
  MUX2IX1 U72 ( .D0(n337), .D1(pmem_twlb[1]), .S(n36), .Y(n34) );
  OAI21BBX1 U73 ( .A(n335), .B(n338), .C(n35), .Y(n646) );
  MUX2IXL U74 ( .D0(n337), .D1(pmem_twlb[0]), .S(n36), .Y(n35) );
  INVX1 U75 ( .A(n322), .Y(n385) );
  NAND21X1 U76 ( .B(n357), .A(n315), .Y(n343) );
  NAND21X1 U77 ( .B(n376), .A(n66), .Y(n315) );
  NAND32X1 U78 ( .B(n366), .C(n267), .A(n266), .Y(N853) );
  INVX1 U79 ( .A(n266), .Y(n359) );
  INVX1 U80 ( .A(n377), .Y(n306) );
  AOI21X1 U81 ( .B(n334), .C(we_twlb), .A(N853), .Y(n36) );
  AO21X1 U82 ( .B(n366), .C(n240), .A(n267), .Y(n93) );
  INVX1 U83 ( .A(n379), .Y(n77) );
  INVX1 U84 ( .A(n379), .Y(n76) );
  INVX1 U85 ( .A(n379), .Y(n75) );
  INVX1 U86 ( .A(n379), .Y(n74) );
  INVX1 U87 ( .A(n84), .Y(n73) );
  INVX1 U88 ( .A(n379), .Y(n72) );
  INVX1 U89 ( .A(n379), .Y(n71) );
  INVX1 U90 ( .A(n84), .Y(n70) );
  INVX1 U91 ( .A(n84), .Y(n69) );
  INVX1 U92 ( .A(n379), .Y(n68) );
  INVX1 U93 ( .A(n84), .Y(n67) );
  INVX1 U94 ( .A(n84), .Y(n78) );
  INVX1 U95 ( .A(n84), .Y(n82) );
  INVX1 U96 ( .A(n84), .Y(n81) );
  INVX1 U97 ( .A(n84), .Y(n80) );
  INVX1 U98 ( .A(n84), .Y(n79) );
  INVX1 U99 ( .A(n84), .Y(n83) );
  INVX1 U100 ( .A(n363), .Y(n203) );
  INVX1 U101 ( .A(n282), .Y(n334) );
  INVX1 U102 ( .A(n112), .Y(n239) );
  NAND21X1 U103 ( .B(n321), .A(n334), .Y(n112) );
  INVX1 U104 ( .A(n354), .Y(n325) );
  INVX1 U105 ( .A(n311), .Y(n386) );
  INVX1 U106 ( .A(n268), .Y(n364) );
  NAND21X1 U107 ( .B(n336), .A(n385), .Y(n268) );
  INVX1 U108 ( .A(n323), .Y(n338) );
  NAND21X1 U109 ( .B(n322), .A(n321), .Y(n323) );
  INVX1 U110 ( .A(n376), .Y(n351) );
  NAND21X1 U111 ( .B(n233), .A(n396), .Y(n377) );
  NAND6XL U112 ( .A(n228), .B(n227), .C(n226), .D(n225), .E(n224), .F(n223), 
        .Y(n240) );
  AND4X1 U113 ( .A(n222), .B(n221), .C(n220), .D(n219), .Y(n223) );
  AND4X1 U114 ( .A(n1), .B(n218), .C(n217), .D(n216), .Y(n224) );
  OAI211X1 U115 ( .C(n236), .D(n231), .A(n348), .B(n396), .Y(n349) );
  INVX1 U116 ( .A(n303), .Y(n231) );
  NAND31X1 U117 ( .C(n316), .A(n38), .B(n39), .Y(n267) );
  AOI21X1 U118 ( .B(n313), .C(n394), .A(n239), .Y(n38) );
  NAND2X1 U119 ( .A(n438), .B(n87), .Y(n281) );
  AND2X1 U120 ( .A(n345), .B(n87), .Y(n39) );
  AO21X1 U121 ( .B(n265), .C(n258), .A(n260), .Y(N894) );
  AO21X1 U122 ( .B(n54), .C(n264), .A(n28), .Y(N889) );
  AO21X1 U123 ( .B(n54), .C(n258), .A(n29), .Y(N886) );
  AO21X1 U124 ( .B(n249), .C(n264), .A(n260), .Y(N885) );
  AO21X1 U125 ( .B(n249), .C(n258), .A(n28), .Y(N882) );
  AO21X1 U126 ( .B(n247), .C(n264), .A(n29), .Y(N881) );
  AO21X1 U127 ( .B(n247), .C(n258), .A(n260), .Y(N878) );
  AND4X1 U128 ( .A(n215), .B(n214), .C(n213), .D(n212), .Y(n225) );
  INVX1 U129 ( .A(n382), .Y(n87) );
  INVX1 U130 ( .A(n314), .Y(n357) );
  NAND21X1 U131 ( .B(n376), .A(n313), .Y(n314) );
  INVX1 U132 ( .A(n269), .Y(n263) );
  INVX1 U133 ( .A(n216), .Y(n165) );
  NAND21X1 U134 ( .B(n346), .A(n345), .Y(n358) );
  OAI211X1 U135 ( .C(n734), .D(n377), .A(n370), .B(n388), .Y(n363) );
  INVX1 U136 ( .A(n234), .Y(n366) );
  NAND21X1 U137 ( .B(n233), .A(n346), .Y(n234) );
  NAND21X1 U138 ( .B(n111), .A(n336), .Y(n282) );
  INVX1 U139 ( .A(n262), .Y(n336) );
  NAND32X1 U140 ( .B(n322), .C(n262), .A(n330), .Y(n354) );
  INVX1 U141 ( .A(n237), .Y(n236) );
  OR2X1 U142 ( .A(n726), .B(n382), .Y(n376) );
  INVX1 U143 ( .A(n341), .Y(n318) );
  NAND2X1 U144 ( .A(n735), .B(n736), .Y(n273) );
  INVX1 U145 ( .A(n340), .Y(n342) );
  INVX1 U146 ( .A(srst), .Y(n88) );
  INVX1 U147 ( .A(n330), .Y(n321) );
  INVX1 U148 ( .A(n734), .Y(n307) );
  INVX1 U149 ( .A(n370), .Y(n278) );
  INVX1 U150 ( .A(n361), .Y(n367) );
  INVX1 U151 ( .A(n150), .Y(n179) );
  INVX1 U152 ( .A(n726), .Y(n394) );
  INVX1 U153 ( .A(n111), .Y(n395) );
  INVX1 U154 ( .A(n389), .Y(n346) );
  INVX1 U155 ( .A(n371), .Y(n316) );
  INVX1 U156 ( .A(n736), .Y(n397) );
  INVX1 U157 ( .A(n360), .Y(n398) );
  AO21X1 U158 ( .B(n107), .C(n388), .A(n382), .Y(n108) );
  OR2X1 U159 ( .A(n726), .B(n312), .Y(n345) );
  NAND21X1 U160 ( .B(n411), .A(n61), .Y(n227) );
  OA222X1 U161 ( .A(memaddr_c[11]), .B(n187), .C(n186), .D(n185), .E(
        memaddr_c[10]), .F(n184), .Y(n191) );
  INVX1 U162 ( .A(n214), .Y(n186) );
  NAND21X1 U163 ( .B(n412), .A(n159), .Y(n210) );
  OA22X1 U164 ( .A(memaddr_c[0]), .B(n209), .C(memaddr_c[1]), .D(n159), .Y(
        n161) );
  INVX1 U165 ( .A(n212), .Y(n194) );
  NAND21X1 U166 ( .B(n191), .A(n215), .Y(n193) );
  NAND32X1 U167 ( .B(n161), .C(n160), .A(n210), .Y(n162) );
  AO21X1 U168 ( .B(N432), .C(n359), .A(n347), .Y(N827) );
  AO21XL U169 ( .B(n358), .C(memaddr_c[1]), .A(n85), .Y(n347) );
  OAI21BBX1 U170 ( .A(N433), .B(n20), .C(n41), .Y(N828) );
  AOI21XL U171 ( .B(n16), .C(memaddr_c[2]), .A(n85), .Y(n41) );
  OAI21BBX1 U172 ( .A(N435), .B(n20), .C(n42), .Y(N830) );
  AOI21XL U173 ( .B(n16), .C(memaddr_c[4]), .A(n26), .Y(n42) );
  OAI21BBX1 U174 ( .A(N436), .B(n20), .C(n43), .Y(N831) );
  AOI21XL U175 ( .B(n16), .C(memaddr_c[5]), .A(n27), .Y(n43) );
  OAI21BBX1 U176 ( .A(N437), .B(n20), .C(n44), .Y(N832) );
  OAI21BBX1 U177 ( .A(N438), .B(n359), .C(n45), .Y(N833) );
  AOI21X1 U178 ( .B(n358), .C(memaddr_c[7]), .A(n27), .Y(n45) );
  OAI21BBX1 U179 ( .A(N441), .B(n359), .C(n46), .Y(N836) );
  AOI21X1 U180 ( .B(n358), .C(memaddr_c[10]), .A(n85), .Y(n46) );
  OAI21BBX1 U181 ( .A(N442), .B(n359), .C(n47), .Y(N837) );
  AOI21X1 U182 ( .B(n358), .C(memaddr_c[11]), .A(n26), .Y(n47) );
  OAI21BBX1 U183 ( .A(N443), .B(n359), .C(n48), .Y(N838) );
  AOI21X1 U184 ( .B(n358), .C(memaddr_c[12]), .A(n27), .Y(n48) );
  OAI21BBX1 U185 ( .A(N444), .B(n359), .C(n49), .Y(N839) );
  AOI21X1 U186 ( .B(n358), .C(memaddr_c[13]), .A(n85), .Y(n49) );
  OAI21BBX1 U187 ( .A(N440), .B(n359), .C(n50), .Y(N835) );
  AOI21X1 U188 ( .B(n358), .C(memaddr_c[9]), .A(n26), .Y(n50) );
  OAI21BBX1 U189 ( .A(N439), .B(n359), .C(n51), .Y(N834) );
  AOI21X1 U190 ( .B(n358), .C(memaddr_c[8]), .A(n27), .Y(n51) );
  OAI21BBX1 U191 ( .A(N434), .B(n20), .C(n52), .Y(N829) );
  AOI21XL U192 ( .B(n16), .C(memaddr_c[3]), .A(n85), .Y(n52) );
  AO21X1 U193 ( .B(n261), .C(n265), .A(n28), .Y(N896) );
  AO21X1 U194 ( .B(n259), .C(n265), .A(n29), .Y(N895) );
  AO21X1 U195 ( .B(n255), .C(n264), .A(n260), .Y(N893) );
  AO21X1 U196 ( .B(n255), .C(n261), .A(n28), .Y(N892) );
  AO21X1 U197 ( .B(n255), .C(n259), .A(n29), .Y(N891) );
  AO21X1 U198 ( .B(n255), .C(n258), .A(n260), .Y(N890) );
  AO21X1 U199 ( .B(n54), .C(n261), .A(n28), .Y(N888) );
  AO21X1 U200 ( .B(n54), .C(n259), .A(n29), .Y(N887) );
  AO21X1 U201 ( .B(n249), .C(n261), .A(n260), .Y(N884) );
  AO21X1 U202 ( .B(n249), .C(n259), .A(n28), .Y(N883) );
  AO21X1 U203 ( .B(n247), .C(n261), .A(n29), .Y(N880) );
  AO21X1 U204 ( .B(n247), .C(n259), .A(n260), .Y(N879) );
  AO21X1 U205 ( .B(n245), .C(n264), .A(n28), .Y(N877) );
  AO21X1 U206 ( .B(n245), .C(n261), .A(n29), .Y(N876) );
  AO21X1 U207 ( .B(n245), .C(n259), .A(n260), .Y(N875) );
  AO21X1 U208 ( .B(n245), .C(n258), .A(n28), .Y(N874) );
  NAND31X1 U209 ( .C(n359), .A(n53), .B(n39), .Y(N825) );
  NAND3XL U210 ( .A(n366), .B(n415), .C(n240), .Y(n53) );
  INVX1 U211 ( .A(n241), .Y(n313) );
  INVX1 U212 ( .A(n217), .Y(n169) );
  INVX1 U213 ( .A(n221), .Y(n171) );
  AOI32XL U214 ( .A(n222), .B(n177), .C(n219), .D(n176), .E(n405), .Y(n183) );
  INVX1 U215 ( .A(n175), .Y(n176) );
  AO21X1 U216 ( .B(n173), .C(n406), .A(n172), .Y(n177) );
  INVX1 U217 ( .A(n174), .Y(n173) );
  INVXL U218 ( .A(memaddr_c[2]), .Y(n411) );
  NAND21X1 U219 ( .B(n410), .A(n63), .Y(n216) );
  NAND21X1 U220 ( .B(n409), .A(n62), .Y(n218) );
  INVX1 U221 ( .A(n292), .Y(n300) );
  NAND21X1 U222 ( .B(n380), .A(n291), .Y(n292) );
  INVX1 U223 ( .A(n285), .Y(n294) );
  NAND21X1 U224 ( .B(n380), .A(n773), .Y(n285) );
  INVX1 U225 ( .A(n286), .Y(n295) );
  NAND21X1 U226 ( .B(n380), .A(n771), .Y(n286) );
  INVX1 U227 ( .A(n287), .Y(n296) );
  NAND21X1 U228 ( .B(n380), .A(n769), .Y(n287) );
  INVX1 U229 ( .A(n289), .Y(n298) );
  NAND21X1 U230 ( .B(n380), .A(n765), .Y(n289) );
  INVX1 U231 ( .A(n290), .Y(n299) );
  NAND21X1 U232 ( .B(n380), .A(n763), .Y(n290) );
  INVX1 U233 ( .A(n284), .Y(n293) );
  NAND21X1 U234 ( .B(n380), .A(n775), .Y(n284) );
  INVX1 U235 ( .A(n288), .Y(n297) );
  NAND21X1 U236 ( .B(n380), .A(n767), .Y(n288) );
  INVX1 U237 ( .A(n252), .Y(n380) );
  INVX1 U238 ( .A(n248), .Y(n249) );
  NAND32X1 U239 ( .B(n251), .C(n250), .A(n373), .Y(n248) );
  INVX1 U240 ( .A(n246), .Y(n247) );
  NAND32X1 U241 ( .B(n373), .C(n250), .A(n251), .Y(n246) );
  NOR3XL U242 ( .A(n373), .B(n251), .C(n250), .Y(n54) );
  INVX1 U243 ( .A(n257), .Y(n265) );
  NAND21X1 U244 ( .B(n373), .A(n256), .Y(n257) );
  INVXL U245 ( .A(memaddr_c[4]), .Y(n409) );
  INVX1 U246 ( .A(memaddr_c[8]), .Y(n405) );
  NAND21X1 U247 ( .B(n408), .A(n64), .Y(n221) );
  NAND21X1 U248 ( .B(n407), .A(n168), .Y(n217) );
  INVX1 U249 ( .A(memaddr_c[7]), .Y(n406) );
  INVXL U250 ( .A(memaddr_c[5]), .Y(n408) );
  OR2X1 U251 ( .A(memaddr_c[9]), .B(n178), .Y(n182) );
  NAND43X1 U252 ( .B(n394), .C(n239), .D(n205), .A(n204), .Y(N820) );
  AO21X1 U253 ( .B(n746), .C(n397), .A(n752), .Y(n205) );
  AND4X1 U254 ( .A(n386), .B(n398), .C(n203), .D(n389), .Y(n204) );
  NAND21X1 U255 ( .B(n405), .A(n175), .Y(n222) );
  NAND21X1 U256 ( .B(n406), .A(n174), .Y(n219) );
  AND2X1 U257 ( .A(n357), .B(n356), .Y(N842) );
  AND2X1 U258 ( .A(N451), .B(n357), .Y(N845) );
  AND2X1 U259 ( .A(N450), .B(n357), .Y(N844) );
  AND2X1 U260 ( .A(N449), .B(n357), .Y(N843) );
  OAI32X1 U261 ( .A(n305), .B(n710), .C(n307), .D(n304), .E(n384), .Y(n648) );
  NAND32X1 U262 ( .B(n394), .C(n26), .A(n735), .Y(n305) );
  OA21XL U263 ( .B(n391), .C(n303), .A(n302), .Y(n304) );
  GEN2XL U264 ( .D(n734), .E(n735), .C(n26), .B(n391), .A(n374), .Y(n302) );
  INVX1 U265 ( .A(memaddr_c[9]), .Y(n404) );
  NAND21X1 U266 ( .B(n404), .A(n178), .Y(n214) );
  NAND21X1 U267 ( .B(n403), .A(n184), .Y(n220) );
  INVX1 U268 ( .A(memaddr_c[10]), .Y(n403) );
  AO21X1 U269 ( .B(sfr_psr), .C(n110), .A(n396), .Y(n262) );
  INVX1 U270 ( .A(n753), .Y(n110) );
  NAND21X1 U271 ( .B(n402), .A(n187), .Y(n212) );
  NAND21X1 U272 ( .B(n401), .A(n192), .Y(n215) );
  INVX1 U273 ( .A(memaddr_c[14]), .Y(n399) );
  INVX1 U274 ( .A(memaddr_c[11]), .Y(n402) );
  INVX1 U275 ( .A(memaddr_c[13]), .Y(n400) );
  INVX1 U276 ( .A(memaddr_c[12]), .Y(n401) );
  INVX1 U277 ( .A(n138), .Y(n114) );
  INVX1 U278 ( .A(n195), .Y(n196) );
  INVX1 U279 ( .A(n384), .Y(n396) );
  NAND32X1 U280 ( .B(n208), .C(n207), .A(n206), .Y(n237) );
  OR4X1 U281 ( .A(n791), .B(n792), .C(n789), .D(n790), .Y(n208) );
  OR4X1 U282 ( .A(n788), .B(N232), .C(n786), .D(n787), .Y(n207) );
  NOR8XL U283 ( .A(n797), .B(n798), .C(n799), .D(n800), .E(n793), .F(n794), 
        .G(n795), .H(n796), .Y(n206) );
  NAND21X1 U284 ( .B(memaddr_c[14]), .A(n2), .Y(n228) );
  AO21X1 U285 ( .B(n325), .C(n414), .A(n37), .Y(n327) );
  OR3XL U286 ( .A(n325), .B(n364), .C(n55), .Y(N898) );
  AOI21X1 U287 ( .B(n361), .C(n749), .A(n269), .Y(n55) );
  NAND32X1 U288 ( .B(n202), .C(n200), .A(n229), .Y(n438) );
  NAND21X1 U289 ( .B(n414), .A(n385), .Y(n340) );
  INVX1 U290 ( .A(n324), .Y(n328) );
  MUX2AXL U291 ( .D0(n438), .D1(sfr_psr), .S(n415), .Y(sfr_psrack) );
  AO21X1 U292 ( .B(n385), .C(n414), .A(n37), .Y(n341) );
  NAND21X1 U293 ( .B(n751), .A(n86), .Y(n269) );
  AOI21X1 U294 ( .B(n271), .C(n270), .A(n27), .Y(N899) );
  AO21X1 U295 ( .B(n416), .C(n414), .A(n398), .Y(n270) );
  NAND21X1 U296 ( .B(n746), .A(n397), .Y(n271) );
  OR3XL U297 ( .A(n94), .B(n92), .C(n97), .Y(n735) );
  OR2X1 U298 ( .A(n106), .B(n90), .Y(n736) );
  OAI31XL U299 ( .A(n728), .B(n753), .C(n109), .D(n754), .Y(n330) );
  INVX1 U300 ( .A(sfr_psw), .Y(n109) );
  INVX1 U301 ( .A(n759), .Y(n106) );
  AO21X1 U302 ( .B(n86), .C(n393), .A(n392), .Y(N821) );
  NAND32X1 U303 ( .B(n390), .C(n750), .A(n389), .Y(n393) );
  INVX1 U304 ( .A(n391), .Y(n392) );
  INVX1 U305 ( .A(n388), .Y(n390) );
  NAND21X1 U306 ( .B(n92), .A(n91), .Y(n734) );
  OR2X1 U307 ( .A(n90), .B(n201), .Y(n361) );
  NAND32X1 U308 ( .B(n229), .C(n201), .A(n200), .Y(n370) );
  NAND32X1 U309 ( .B(n229), .C(n106), .A(n200), .Y(n388) );
  INVX1 U310 ( .A(n154), .Y(n151) );
  NAND32X1 U311 ( .B(n144), .C(n152), .A(n151), .Y(n150) );
  NAND32X1 U312 ( .B(n146), .C(n189), .A(n188), .Y(n148) );
  INVX1 U313 ( .A(n149), .Y(n188) );
  INVX1 U314 ( .A(n209), .Y(n211) );
  AND4X1 U315 ( .A(n258), .B(n372), .C(n251), .D(n373), .Y(n197) );
  INVX1 U316 ( .A(n238), .Y(n348) );
  INVX1 U317 ( .A(n230), .Y(n258) );
  NAND21X1 U318 ( .B(n97), .A(n759), .Y(n111) );
  OR2X1 U319 ( .A(n229), .B(n276), .Y(n389) );
  AO21X1 U320 ( .B(n201), .C(n202), .A(n97), .Y(n726) );
  NAND21X1 U321 ( .B(n415), .A(n346), .Y(n371) );
  INVX1 U322 ( .A(n275), .Y(n105) );
  INVX1 U323 ( .A(n95), .Y(n103) );
  NAND21X1 U324 ( .B(n279), .A(n105), .Y(n95) );
  INVX1 U325 ( .A(n279), .Y(n104) );
  NAND21X1 U326 ( .B(n367), .A(n107), .Y(n360) );
  NAND21X1 U327 ( .B(n111), .A(n414), .Y(n747) );
  INVX1 U328 ( .A(n749), .Y(n424) );
  INVX1 U329 ( .A(n751), .Y(n368) );
  INVX1 U330 ( .A(n375), .Y(n264) );
  NAND31X1 U331 ( .C(d_psrd), .A(n56), .B(n238), .Y(n241) );
  NAND3XL U332 ( .A(n306), .B(n240), .C(n237), .Y(n56) );
  NAND43X1 U333 ( .B(n236), .C(n235), .D(d_psrd), .A(n306), .Y(n312) );
  INVXL U334 ( .A(n240), .Y(n235) );
  GEN2XL U335 ( .D(c_adr[14]), .E(n399), .C(n141), .B(n140), .A(n139), .Y(n199) );
  AOI21XL U336 ( .B(n228), .C(n213), .A(n197), .Y(n198) );
  OAI32X1 U337 ( .A(n114), .B(memaddr_c[12]), .C(n146), .D(memaddr_c[13]), .E(
        n113), .Y(n141) );
  AO2222XL U338 ( .A(n344), .B(memaddr_c[8]), .C(pre_1_adr[8]), .D(n4), .E(
        memaddr[8]), .F(n342), .G(sfr_psofs[8]), .H(n341), .Y(N862) );
  AO2222XL U339 ( .A(n344), .B(memaddr_c[9]), .C(pre_1_adr[9]), .D(n4), .E(
        memaddr[9]), .F(n342), .G(sfr_psofs[9]), .H(n341), .Y(N863) );
  AND3X1 U340 ( .A(n138), .B(n140), .C(n137), .Y(n139) );
  OA21X1 U341 ( .B(c_adr[12]), .C(n401), .A(n136), .Y(n137) );
  AO21X1 U342 ( .B(c_adr[11]), .C(n402), .A(n135), .Y(n136) );
  GEN2XL U343 ( .D(c_adr[9]), .E(n404), .C(n134), .B(n133), .A(n132), .Y(n135)
         );
  AND3X1 U344 ( .A(pmem_clk[0]), .B(n40), .C(n276), .Y(n274) );
  AO2222XL U345 ( .A(n344), .B(memaddr_c[7]), .C(pre_1_adr[7]), .D(n343), .E(
        memaddr[7]), .F(n342), .G(sfr_psofs[7]), .H(n341), .Y(N861) );
  AO2222XL U346 ( .A(n344), .B(memaddr_c[10]), .C(pre_1_adr[10]), .D(n4), .E(
        memaddr[10]), .F(n342), .G(sfr_psofs[10]), .H(n341), .Y(N864) );
  AO2222XL U347 ( .A(n344), .B(memaddr_c[1]), .C(pre_1_adr[1]), .D(n343), .E(
        memaddr[1]), .F(n342), .G(sfr_psofs[1]), .H(n341), .Y(N855) );
  AO2222XL U348 ( .A(n344), .B(memaddr_c[13]), .C(pre_1_adr[13]), .D(n4), .E(
        memaddr[13]), .F(n342), .G(sfr_psofs[13]), .H(n341), .Y(N867) );
  AO2222XL U349 ( .A(n344), .B(memaddr_c[12]), .C(pre_1_adr[12]), .D(n4), .E(
        memaddr[12]), .F(n342), .G(sfr_psofs[12]), .H(n341), .Y(N866) );
  AO2222XL U350 ( .A(n344), .B(memaddr_c[11]), .C(pre_1_adr[11]), .D(n343), 
        .E(memaddr[11]), .F(n342), .G(sfr_psofs[11]), .H(n341), .Y(N865) );
  AO2222XL U351 ( .A(n21), .B(memaddr_c[6]), .C(pre_1_adr[6]), .D(n4), .E(
        memaddr[6]), .F(n342), .G(sfr_psofs[6]), .H(n341), .Y(N860) );
  AO2222XL U352 ( .A(n21), .B(memaddr_c[5]), .C(pre_1_adr[5]), .D(n343), .E(
        memaddr[5]), .F(n342), .G(sfr_psofs[5]), .H(n24), .Y(N859) );
  AO2222XL U353 ( .A(n21), .B(memaddr_c[4]), .C(pre_1_adr[4]), .D(n4), .E(
        memaddr[4]), .F(n15), .G(sfr_psofs[4]), .H(n24), .Y(N858) );
  AO2222XL U354 ( .A(n21), .B(memaddr_c[3]), .C(pre_1_adr[3]), .D(n343), .E(
        memaddr[3]), .F(n15), .G(sfr_psofs[3]), .H(n24), .Y(N857) );
  AO2222XL U355 ( .A(n21), .B(memaddr_c[2]), .C(pre_1_adr[2]), .D(n4), .E(
        memaddr[2]), .F(n15), .G(sfr_psofs[2]), .H(n24), .Y(N856) );
  AO2222XL U356 ( .A(n21), .B(memaddr_c[0]), .C(pre_1_adr[0]), .D(n343), .E(
        memaddr[0]), .F(n15), .G(sfr_psofs[0]), .H(n24), .Y(N854) );
  AND3X1 U357 ( .A(wd_twlb[0]), .B(we_twlb), .C(n336), .Y(n335) );
  AND3X1 U358 ( .A(wd_twlb[1]), .B(we_twlb), .C(n336), .Y(n339) );
  OAI21BBX1 U359 ( .A(N445), .B(n359), .C(n57), .Y(N840) );
  AOI21X1 U360 ( .B(n358), .C(memaddr_c[14]), .A(n85), .Y(n57) );
  OAI21BBX1 U361 ( .A(N431), .B(n20), .C(n58), .Y(N826) );
  INVX1 U362 ( .A(n435), .Y(n118) );
  OAI32X1 U363 ( .A(n130), .B(memaddr_c[8]), .C(n144), .D(n129), .E(n128), .Y(
        n134) );
  AO21X1 U364 ( .B(memaddr_c[8]), .C(n144), .A(n130), .Y(n128) );
  AOI211X1 U365 ( .C(c_adr[7]), .D(n406), .A(n127), .B(n126), .Y(n129) );
  INVX1 U366 ( .A(n115), .Y(n130) );
  OAI211X1 U367 ( .C(pre_1_adr[13]), .D(n333), .A(n332), .B(n331), .Y(n337) );
  AOI33X1 U368 ( .A(n330), .B(n329), .C(n328), .D(sfr_psofs[14]), .E(n327), 
        .F(n326), .Y(n331) );
  NAND32X1 U369 ( .B(memaddr_c[13]), .C(n399), .A(n344), .Y(n332) );
  INVX1 U370 ( .A(sfr_psofs[13]), .Y(n326) );
  AOI221XL U371 ( .A(memaddr_c[4]), .B(n432), .C(n125), .D(n124), .E(n123), 
        .Y(n126) );
  AO21XL U372 ( .B(memaddr_c[2]), .C(n119), .A(n118), .Y(n124) );
  INVX1 U373 ( .A(n122), .Y(n125) );
  OAI22AXL U374 ( .D(c_adr[0]), .C(n59), .A(memaddr_c[1]), .B(n430), .Y(n437)
         );
  AO21XL U375 ( .B(memaddr_c[1]), .C(n430), .A(memaddr_c[0]), .Y(n59) );
  OAI211XL U376 ( .C(n399), .D(n320), .A(n333), .B(n319), .Y(N868) );
  OA21X1 U377 ( .B(n318), .C(n317), .A(n324), .Y(n319) );
  INVX1 U378 ( .A(n344), .Y(n320) );
  INVX1 U379 ( .A(sfr_psofs[14]), .Y(n317) );
  NAND21X1 U380 ( .B(d_psrd), .A(n241), .Y(n252) );
  NAND32X1 U381 ( .B(c_ptr[4]), .C(n376), .A(n252), .Y(n250) );
  INVX1 U382 ( .A(n434), .Y(n117) );
  AO21X1 U383 ( .B(dbg_01[0]), .C(n83), .A(n30), .Y(N479) );
  AO21X1 U384 ( .B(dbg_02[0]), .C(n83), .A(n31), .Y(N487) );
  AO21X1 U385 ( .B(dbg_03[0]), .C(n83), .A(n293), .Y(N495) );
  AO21X1 U386 ( .B(dbg_04[0]), .C(n83), .A(n30), .Y(N503) );
  AO21X1 U387 ( .B(dbg_05[0]), .C(n83), .A(n31), .Y(N511) );
  AO21X1 U388 ( .B(dbg_06[0]), .C(n83), .A(n293), .Y(N519) );
  AO21X1 U389 ( .B(n78), .C(dbg_07[0]), .A(n30), .Y(N527) );
  AO21X1 U390 ( .B(dbg_01[1]), .C(n82), .A(n22), .Y(N480) );
  AO21X1 U391 ( .B(dbg_02[1]), .C(n82), .A(n23), .Y(N488) );
  AO21X1 U392 ( .B(dbg_03[1]), .C(n82), .A(n294), .Y(N496) );
  AO21X1 U393 ( .B(dbg_04[1]), .C(n82), .A(n22), .Y(N504) );
  AO21X1 U394 ( .B(dbg_05[1]), .C(n82), .A(n23), .Y(N512) );
  AO21X1 U395 ( .B(dbg_06[1]), .C(n82), .A(n294), .Y(N520) );
  AO21X1 U396 ( .B(n78), .C(dbg_07[1]), .A(n22), .Y(N528) );
  AO21X1 U397 ( .B(dbg_01[2]), .C(n82), .A(n17), .Y(N481) );
  AO21X1 U398 ( .B(dbg_02[2]), .C(n82), .A(n18), .Y(N489) );
  AO21X1 U399 ( .B(dbg_03[2]), .C(n82), .A(n295), .Y(N497) );
  AO21X1 U400 ( .B(dbg_04[2]), .C(n81), .A(n17), .Y(N505) );
  AO21X1 U401 ( .B(dbg_05[2]), .C(n82), .A(n18), .Y(N513) );
  AO21X1 U402 ( .B(dbg_06[2]), .C(n81), .A(n295), .Y(N521) );
  AO21X1 U403 ( .B(n78), .C(dbg_07[2]), .A(n17), .Y(N529) );
  AO21X1 U404 ( .B(dbg_01[3]), .C(n81), .A(n13), .Y(N482) );
  AO21X1 U405 ( .B(dbg_02[3]), .C(n81), .A(n14), .Y(N490) );
  AO21X1 U406 ( .B(dbg_03[3]), .C(n81), .A(n296), .Y(N498) );
  AO21X1 U407 ( .B(dbg_04[3]), .C(n81), .A(n13), .Y(N506) );
  AO21X1 U408 ( .B(dbg_05[3]), .C(n81), .A(n14), .Y(N514) );
  AO21X1 U409 ( .B(dbg_06[3]), .C(n81), .A(n296), .Y(N522) );
  AO21X1 U410 ( .B(n78), .C(dbg_07[3]), .A(n13), .Y(N530) );
  AO21X1 U411 ( .B(dbg_01[4]), .C(n80), .A(n11), .Y(N483) );
  AO21X1 U412 ( .B(dbg_02[4]), .C(n80), .A(n12), .Y(N491) );
  AO21X1 U413 ( .B(dbg_03[4]), .C(n81), .A(n297), .Y(N499) );
  AO21X1 U414 ( .B(dbg_04[4]), .C(n80), .A(n11), .Y(N507) );
  AO21X1 U415 ( .B(dbg_05[4]), .C(n80), .A(n12), .Y(N515) );
  AO21X1 U416 ( .B(dbg_06[4]), .C(n81), .A(n297), .Y(N523) );
  AO21X1 U417 ( .B(n78), .C(dbg_07[4]), .A(n11), .Y(N531) );
  AO21X1 U418 ( .B(dbg_01[5]), .C(n80), .A(n9), .Y(N484) );
  AO21X1 U419 ( .B(dbg_02[5]), .C(n80), .A(n10), .Y(N492) );
  AO21X1 U420 ( .B(dbg_03[5]), .C(n80), .A(n298), .Y(N500) );
  AO21X1 U421 ( .B(dbg_04[5]), .C(n80), .A(n9), .Y(N508) );
  AO21X1 U422 ( .B(dbg_05[5]), .C(n80), .A(n10), .Y(N516) );
  AO21X1 U423 ( .B(dbg_06[5]), .C(n79), .A(n298), .Y(N524) );
  AO21X1 U424 ( .B(n78), .C(dbg_07[5]), .A(n9), .Y(N532) );
  AO21X1 U425 ( .B(dbg_01[6]), .C(n80), .A(n7), .Y(N485) );
  AO21X1 U426 ( .B(dbg_02[6]), .C(n79), .A(n8), .Y(N493) );
  AO21X1 U427 ( .B(dbg_03[6]), .C(n79), .A(n299), .Y(N501) );
  AO21X1 U428 ( .B(dbg_04[6]), .C(n79), .A(n7), .Y(N509) );
  AO21X1 U429 ( .B(dbg_05[6]), .C(n79), .A(n8), .Y(N517) );
  AO21X1 U430 ( .B(dbg_06[6]), .C(n79), .A(n299), .Y(N525) );
  AO21X1 U431 ( .B(n78), .C(dbg_07[6]), .A(n7), .Y(N533) );
  AO21X1 U432 ( .B(dbg_01[7]), .C(n79), .A(n5), .Y(N486) );
  AO21X1 U433 ( .B(dbg_02[7]), .C(n79), .A(n6), .Y(N494) );
  AO21X1 U434 ( .B(dbg_03[7]), .C(n79), .A(n300), .Y(N502) );
  AO21X1 U435 ( .B(dbg_04[7]), .C(n78), .A(n5), .Y(N510) );
  AO21X1 U436 ( .B(dbg_05[7]), .C(n78), .A(n6), .Y(N518) );
  AO21X1 U437 ( .B(dbg_06[7]), .C(n79), .A(n300), .Y(N526) );
  AO21X1 U438 ( .B(n78), .C(dbg_07[7]), .A(n5), .Y(N534) );
  AO21X1 U439 ( .B(n77), .C(dbg_08[0]), .A(n31), .Y(N535) );
  AO21X1 U440 ( .B(n77), .C(dbg_08[1]), .A(n23), .Y(N536) );
  AO21X1 U441 ( .B(n77), .C(dbg_08[2]), .A(n18), .Y(N537) );
  AO21X1 U442 ( .B(n77), .C(dbg_08[3]), .A(n14), .Y(N538) );
  AO21X1 U443 ( .B(n77), .C(dbg_08[4]), .A(n12), .Y(N539) );
  AO21X1 U444 ( .B(n77), .C(dbg_08[5]), .A(n10), .Y(N540) );
  AO21X1 U445 ( .B(n77), .C(dbg_08[6]), .A(n8), .Y(N541) );
  AO21X1 U446 ( .B(n77), .C(dbg_08[7]), .A(n6), .Y(N542) );
  AO21X1 U447 ( .B(n77), .C(dbg_09[0]), .A(n293), .Y(N543) );
  AO21X1 U448 ( .B(n77), .C(dbg_09[1]), .A(n294), .Y(N544) );
  AO21X1 U449 ( .B(n76), .C(dbg_09[2]), .A(n295), .Y(N545) );
  AO21X1 U450 ( .B(n76), .C(dbg_09[3]), .A(n296), .Y(N546) );
  AO21X1 U451 ( .B(n76), .C(dbg_09[4]), .A(n297), .Y(N547) );
  AO21X1 U452 ( .B(n76), .C(dbg_09[5]), .A(n298), .Y(N548) );
  AO21X1 U453 ( .B(n76), .C(dbg_09[6]), .A(n299), .Y(N549) );
  AO21X1 U454 ( .B(n76), .C(dbg_09[7]), .A(n300), .Y(N550) );
  AO21X1 U455 ( .B(n76), .C(dbg_0a[0]), .A(n30), .Y(N551) );
  AO21X1 U456 ( .B(n76), .C(dbg_0a[1]), .A(n22), .Y(N552) );
  AO21X1 U457 ( .B(n76), .C(dbg_0a[2]), .A(n17), .Y(N553) );
  AO21X1 U458 ( .B(n76), .C(dbg_0a[3]), .A(n13), .Y(N554) );
  AO21X1 U459 ( .B(n75), .C(dbg_0a[4]), .A(n11), .Y(N555) );
  AO21X1 U460 ( .B(n75), .C(dbg_0a[5]), .A(n9), .Y(N556) );
  AO21X1 U461 ( .B(n75), .C(dbg_0a[6]), .A(n7), .Y(N557) );
  AO21X1 U462 ( .B(n75), .C(dbg_0a[7]), .A(n5), .Y(N558) );
  AO21X1 U463 ( .B(n75), .C(dbg_0b[0]), .A(n31), .Y(N559) );
  AO21X1 U464 ( .B(n75), .C(dbg_0b[1]), .A(n23), .Y(N560) );
  AO21X1 U465 ( .B(n75), .C(dbg_0b[2]), .A(n18), .Y(N561) );
  AO21X1 U466 ( .B(n75), .C(dbg_0b[3]), .A(n14), .Y(N562) );
  AO21X1 U467 ( .B(n75), .C(dbg_0b[4]), .A(n12), .Y(N563) );
  AO21X1 U468 ( .B(n75), .C(dbg_0b[5]), .A(n10), .Y(N564) );
  AO21X1 U469 ( .B(n301), .C(dbg_0b[6]), .A(n8), .Y(N565) );
  AO21X1 U470 ( .B(n301), .C(dbg_0b[7]), .A(n6), .Y(N566) );
  AO21X1 U471 ( .B(n83), .C(dbg_0c[0]), .A(n293), .Y(N567) );
  AO21X1 U472 ( .B(n83), .C(dbg_0c[1]), .A(n294), .Y(N568) );
  AO21X1 U473 ( .B(n301), .C(dbg_0c[2]), .A(n295), .Y(N569) );
  AO21X1 U474 ( .B(n301), .C(dbg_0c[3]), .A(n296), .Y(N570) );
  AO21X1 U475 ( .B(n83), .C(dbg_0c[4]), .A(n297), .Y(N571) );
  AO21X1 U476 ( .B(n301), .C(dbg_0c[5]), .A(n298), .Y(N572) );
  AO21X1 U477 ( .B(n301), .C(dbg_0c[6]), .A(n299), .Y(N573) );
  AO21X1 U478 ( .B(n74), .C(dbg_0c[7]), .A(n300), .Y(N574) );
  AO21X1 U479 ( .B(n74), .C(dbg_0d[0]), .A(n30), .Y(N575) );
  AO21X1 U480 ( .B(n74), .C(dbg_0d[1]), .A(n22), .Y(N576) );
  AO21X1 U481 ( .B(n74), .C(dbg_0d[2]), .A(n17), .Y(N577) );
  AO21X1 U482 ( .B(n74), .C(dbg_0d[3]), .A(n13), .Y(N578) );
  AO21X1 U483 ( .B(n74), .C(dbg_0d[4]), .A(n11), .Y(N579) );
  AO21X1 U484 ( .B(n74), .C(dbg_0d[5]), .A(n9), .Y(N580) );
  AO21X1 U485 ( .B(n74), .C(dbg_0d[6]), .A(n7), .Y(N581) );
  AO21X1 U486 ( .B(n74), .C(dbg_0d[7]), .A(n5), .Y(N582) );
  AO21X1 U487 ( .B(n74), .C(dbg_0e[0]), .A(n31), .Y(N583) );
  AO21X1 U488 ( .B(n73), .C(dbg_0e[1]), .A(n23), .Y(N584) );
  AO21X1 U489 ( .B(n73), .C(dbg_0e[2]), .A(n18), .Y(N585) );
  AO21X1 U490 ( .B(n73), .C(dbg_0e[3]), .A(n14), .Y(N586) );
  AO21X1 U491 ( .B(n73), .C(dbg_0e[4]), .A(n12), .Y(N587) );
  AO21X1 U492 ( .B(n73), .C(dbg_0e[5]), .A(n10), .Y(N588) );
  AO21X1 U493 ( .B(n73), .C(dbg_0e[6]), .A(n8), .Y(N589) );
  AO21X1 U494 ( .B(n73), .C(dbg_0e[7]), .A(n6), .Y(N590) );
  AO21X1 U495 ( .B(n73), .C(dbg_0f[0]), .A(n293), .Y(N591) );
  AO21X1 U496 ( .B(n73), .C(dbg_0f[1]), .A(n294), .Y(N592) );
  AO21X1 U497 ( .B(n73), .C(dbg_0f[2]), .A(n295), .Y(N593) );
  AO21X1 U498 ( .B(n72), .C(dbg_0f[3]), .A(n296), .Y(N594) );
  AO21X1 U499 ( .B(n72), .C(dbg_0f[4]), .A(n297), .Y(N595) );
  AO21X1 U500 ( .B(n72), .C(dbg_0f[5]), .A(n298), .Y(N596) );
  AO21X1 U501 ( .B(n72), .C(dbg_0f[6]), .A(n299), .Y(N597) );
  AO21X1 U502 ( .B(n72), .C(dbg_0f[7]), .A(n300), .Y(N598) );
  AO21X1 U503 ( .B(n72), .C(c_buf_16__0_), .A(n30), .Y(N599) );
  AO21X1 U504 ( .B(n72), .C(c_buf_16__1_), .A(n22), .Y(N600) );
  AO21X1 U505 ( .B(n72), .C(c_buf_16__2_), .A(n17), .Y(N601) );
  AO21X1 U506 ( .B(n72), .C(c_buf_16__3_), .A(n13), .Y(N602) );
  AO21X1 U507 ( .B(n72), .C(c_buf_16__4_), .A(n11), .Y(N603) );
  AO21X1 U508 ( .B(n71), .C(c_buf_16__5_), .A(n9), .Y(N604) );
  AO21X1 U509 ( .B(n71), .C(c_buf_16__6_), .A(n7), .Y(N605) );
  AO21X1 U510 ( .B(n71), .C(c_buf_16__7_), .A(n5), .Y(N606) );
  AO21X1 U511 ( .B(n71), .C(c_buf_17__0_), .A(n31), .Y(N607) );
  AO21X1 U512 ( .B(n71), .C(c_buf_17__1_), .A(n23), .Y(N608) );
  AO21X1 U513 ( .B(n71), .C(c_buf_17__2_), .A(n18), .Y(N609) );
  AO21X1 U514 ( .B(n71), .C(c_buf_17__3_), .A(n14), .Y(N610) );
  AO21X1 U515 ( .B(n71), .C(c_buf_17__4_), .A(n12), .Y(N611) );
  AO21X1 U516 ( .B(n71), .C(c_buf_17__5_), .A(n10), .Y(N612) );
  AO21X1 U517 ( .B(n71), .C(c_buf_17__6_), .A(n8), .Y(N613) );
  AO21X1 U518 ( .B(n70), .C(c_buf_17__7_), .A(n6), .Y(N614) );
  AO21X1 U519 ( .B(n70), .C(c_buf_18__0_), .A(n293), .Y(N615) );
  AO21X1 U520 ( .B(n70), .C(c_buf_18__1_), .A(n294), .Y(N616) );
  AO21X1 U521 ( .B(n70), .C(c_buf_18__2_), .A(n295), .Y(N617) );
  AO21X1 U522 ( .B(n70), .C(c_buf_18__3_), .A(n296), .Y(N618) );
  AO21X1 U523 ( .B(n70), .C(c_buf_18__4_), .A(n297), .Y(N619) );
  AO21X1 U524 ( .B(n70), .C(c_buf_18__5_), .A(n298), .Y(N620) );
  AO21X1 U525 ( .B(n70), .C(c_buf_18__6_), .A(n299), .Y(N621) );
  AO21X1 U526 ( .B(n70), .C(c_buf_18__7_), .A(n300), .Y(N622) );
  AO21X1 U527 ( .B(n70), .C(c_buf_19__0_), .A(n30), .Y(N623) );
  AO21X1 U528 ( .B(n69), .C(c_buf_19__1_), .A(n22), .Y(N624) );
  AO21X1 U529 ( .B(n69), .C(c_buf_19__2_), .A(n17), .Y(N625) );
  AO21X1 U530 ( .B(n69), .C(c_buf_19__3_), .A(n13), .Y(N626) );
  AO21X1 U531 ( .B(n69), .C(c_buf_19__4_), .A(n11), .Y(N627) );
  AO21X1 U532 ( .B(n69), .C(c_buf_19__5_), .A(n9), .Y(N628) );
  AO21X1 U533 ( .B(n69), .C(c_buf_19__6_), .A(n7), .Y(N629) );
  AO21X1 U534 ( .B(n69), .C(c_buf_19__7_), .A(n5), .Y(N630) );
  AO21X1 U535 ( .B(n69), .C(c_buf_20__0_), .A(n31), .Y(N631) );
  AO21X1 U536 ( .B(n69), .C(c_buf_20__1_), .A(n23), .Y(N632) );
  AO21X1 U537 ( .B(n69), .C(c_buf_20__2_), .A(n18), .Y(N633) );
  AO21X1 U538 ( .B(n68), .C(c_buf_20__3_), .A(n14), .Y(N634) );
  AO21X1 U539 ( .B(n68), .C(c_buf_20__4_), .A(n12), .Y(N635) );
  AO21X1 U540 ( .B(n68), .C(c_buf_20__5_), .A(n10), .Y(N636) );
  AO21X1 U541 ( .B(n68), .C(c_buf_20__6_), .A(n8), .Y(N637) );
  AO21X1 U542 ( .B(n68), .C(c_buf_20__7_), .A(n6), .Y(N638) );
  AO21X1 U543 ( .B(n68), .C(c_buf_21__0_), .A(n293), .Y(N639) );
  AO21X1 U544 ( .B(n68), .C(c_buf_21__1_), .A(n294), .Y(N640) );
  AO21X1 U545 ( .B(n68), .C(c_buf_21__2_), .A(n295), .Y(N641) );
  AO21X1 U546 ( .B(n68), .C(c_buf_21__3_), .A(n296), .Y(N642) );
  AO21X1 U547 ( .B(n68), .C(c_buf_21__4_), .A(n297), .Y(N643) );
  AO21X1 U548 ( .B(n67), .C(c_buf_21__5_), .A(n298), .Y(N644) );
  AO21X1 U549 ( .B(n67), .C(c_buf_21__6_), .A(n299), .Y(N645) );
  AO21X1 U550 ( .B(n67), .C(c_buf_21__7_), .A(n300), .Y(N646) );
  AO21X1 U551 ( .B(n67), .C(c_buf_22__0_), .A(n30), .Y(N647) );
  AO21X1 U552 ( .B(n67), .C(c_buf_22__1_), .A(n22), .Y(N648) );
  AO21X1 U553 ( .B(n67), .C(c_buf_22__2_), .A(n17), .Y(N649) );
  AO21X1 U554 ( .B(n67), .C(c_buf_22__3_), .A(n13), .Y(N650) );
  AO21X1 U555 ( .B(n67), .C(c_buf_22__4_), .A(n11), .Y(N651) );
  AO21X1 U556 ( .B(n67), .C(c_buf_22__5_), .A(n9), .Y(N652) );
  AO21X1 U557 ( .B(n67), .C(c_buf_22__6_), .A(n7), .Y(N653) );
  AO21XL U558 ( .B(n66), .C(c_buf_22__7_), .A(n300), .Y(N654) );
  AO21XL U559 ( .B(n66), .C(wr_buf[0]), .A(n293), .Y(N655) );
  AO21XL U560 ( .B(n66), .C(wr_buf[1]), .A(n294), .Y(N656) );
  AO21XL U561 ( .B(n66), .C(wr_buf[2]), .A(n295), .Y(N657) );
  AO21XL U562 ( .B(n66), .C(wr_buf[3]), .A(n296), .Y(N658) );
  AO21XL U563 ( .B(n66), .C(wr_buf[4]), .A(n297), .Y(N659) );
  AO21XL U564 ( .B(n66), .C(wr_buf[5]), .A(n298), .Y(N660) );
  AO21XL U565 ( .B(n66), .C(wr_buf[6]), .A(n299), .Y(N661) );
  AO21X1 U566 ( .B(n83), .C(wr_buf[7]), .A(n5), .Y(N662) );
  OA21XL U567 ( .B(n748), .C(r_pwdn_en), .A(n349), .Y(n352) );
  NAND21X1 U568 ( .B(n355), .A(n354), .Y(N824) );
  GEN2XL U569 ( .D(n353), .E(n352), .C(n25), .B(n351), .A(n350), .Y(n355) );
  OA21X1 U570 ( .B(n19), .C(n360), .A(n86), .Y(n350) );
  AND3X1 U571 ( .A(n348), .B(cs_ft[0]), .C(n377), .Y(n353) );
  INVX1 U572 ( .A(n253), .Y(n256) );
  NAND43X1 U573 ( .B(c_ptr[3]), .C(n380), .D(n376), .A(c_ptr[4]), .Y(n253) );
  OAI21X1 U574 ( .B(n383), .C(n26), .A(n381), .Y(N822) );
  AND4X1 U575 ( .A(n371), .B(n370), .C(n735), .D(n369), .Y(n383) );
  GEN2XL U576 ( .D(n380), .E(n379), .C(n378), .B(n377), .A(n376), .Y(n381) );
  AOI221XL U577 ( .A(n368), .B(n424), .C(n367), .D(mcu_psw), .E(n366), .Y(n369) );
  INVX1 U578 ( .A(n242), .Y(n245) );
  NAND32X1 U579 ( .B(c_ptr[3]), .C(n250), .A(n373), .Y(n242) );
  INVX1 U580 ( .A(n254), .Y(n255) );
  NAND21X1 U581 ( .B(c_ptr[2]), .A(n256), .Y(n254) );
  AO21X1 U582 ( .B(n86), .C(n365), .A(n364), .Y(N823) );
  NAND32X1 U583 ( .B(n397), .C(n363), .A(n362), .Y(n365) );
  AOI32X1 U584 ( .A(n361), .B(mcu_psw), .C(n360), .D(n368), .E(n749), .Y(n362)
         );
  AND2X1 U585 ( .A(N452), .B(n357), .Y(N846) );
  OAI32XL U586 ( .A(memaddr_c[6]), .B(n143), .C(n117), .D(n116), .E(n120), .Y(
        n127) );
  AOI32X1 U587 ( .A(n436), .B(c_adr[4]), .C(n409), .D(c_adr[5]), .E(n408), .Y(
        n116) );
  NAND21X1 U588 ( .B(c_adr[9]), .A(memaddr_c[9]), .Y(n115) );
  NAND21X1 U589 ( .B(c_adr[11]), .A(memaddr_c[11]), .Y(n131) );
  AO21X1 U590 ( .B(n385), .C(n311), .A(n310), .Y(n647) );
  MUX2BXL U591 ( .D0(n309), .D1(n308), .S(n307), .Y(n310) );
  AND2X1 U592 ( .A(pmem_re), .B(n386), .Y(n309) );
  NAND21X1 U593 ( .B(n27), .A(n306), .Y(n308) );
  OA21X1 U594 ( .B(c_adr[10]), .C(n403), .A(n131), .Y(n133) );
  NOR6XL U595 ( .A(c_ptr[3]), .B(n375), .C(n374), .D(n25), .E(n373), .F(n372), 
        .Y(n378) );
  NAND21X1 U596 ( .B(c_adr[13]), .A(memaddr_c[13]), .Y(n138) );
  NAND2X1 U597 ( .A(hit_ps_c), .B(mcu_psr_c), .Y(n384) );
  AND3X1 U598 ( .A(c_adr[10]), .B(n403), .C(n131), .Y(n132) );
  INVX1 U599 ( .A(cs_n), .Y(pmem_csb) );
  NAND21X1 U600 ( .B(c_adr[14]), .A(memaddr_c[14]), .Y(n140) );
  MUX2X1 U601 ( .D0(pmem_pgm), .D1(n385), .S(n60), .Y(n644) );
  NAND2X1 U602 ( .A(n283), .B(n282), .Y(n60) );
  MUX2X1 U603 ( .D0(n387), .D1(n25), .S(n386), .Y(n649) );
  AND2X1 U604 ( .A(n385), .B(n384), .Y(n387) );
  INVX1 U605 ( .A(dbg_07[7]), .Y(n488) );
  INVX1 U606 ( .A(dbg_08[7]), .Y(n490) );
  INVX1 U607 ( .A(dbg_09[7]), .Y(n492) );
  INVX1 U608 ( .A(c_buf_21__7_), .Y(n459) );
  INVX1 U609 ( .A(c_buf_22__7_), .Y(n461) );
  INVX1 U610 ( .A(c_adr[4]), .Y(n432) );
  INVX1 U611 ( .A(c_adr[3]), .Y(n431) );
  INVX1 U612 ( .A(c_adr[1]), .Y(n430) );
  INVX1 U613 ( .A(c_adr[0]), .Y(n433) );
  INVX1 U614 ( .A(c_buf_21__5_), .Y(n533) );
  INVX1 U615 ( .A(c_buf_22__5_), .Y(n534) );
  INVX1 U616 ( .A(c_buf_21__6_), .Y(n507) );
  INVX1 U617 ( .A(c_buf_22__6_), .Y(n508) );
  INVX1 U618 ( .A(c_buf_21__2_), .Y(n611) );
  INVX1 U619 ( .A(c_buf_22__2_), .Y(n612) );
  INVX1 U620 ( .A(c_buf_21__1_), .Y(n637) );
  INVX1 U621 ( .A(c_buf_22__1_), .Y(n638) );
  INVX1 U622 ( .A(dbg_0a[7]), .Y(n484) );
  INVX1 U623 ( .A(dbg_0b[7]), .Y(n486) );
  INVX1 U624 ( .A(dbg_07[5]), .Y(n548) );
  INVX1 U625 ( .A(dbg_08[5]), .Y(n549) );
  INVX1 U626 ( .A(dbg_09[5]), .Y(n550) );
  INVX1 U627 ( .A(dbg_07[6]), .Y(n522) );
  INVX1 U628 ( .A(dbg_08[6]), .Y(n523) );
  INVX1 U629 ( .A(dbg_09[6]), .Y(n524) );
  INVX1 U630 ( .A(dbg_07[4]), .Y(n574) );
  INVX1 U631 ( .A(dbg_08[4]), .Y(n575) );
  INVX1 U632 ( .A(dbg_09[4]), .Y(n576) );
  INVX1 U633 ( .A(dbg_07[0]), .Y(n698) );
  INVX1 U634 ( .A(dbg_08[0]), .Y(n699) );
  INVX1 U635 ( .A(dbg_09[0]), .Y(n700) );
  INVX1 U636 ( .A(dbg_07[3]), .Y(n600) );
  INVX1 U637 ( .A(dbg_08[3]), .Y(n601) );
  INVX1 U638 ( .A(dbg_09[3]), .Y(n602) );
  INVX1 U639 ( .A(dbg_07[2]), .Y(n626) );
  INVX1 U640 ( .A(dbg_08[2]), .Y(n627) );
  INVX1 U641 ( .A(dbg_09[2]), .Y(n628) );
  INVX1 U642 ( .A(dbg_07[1]), .Y(n663) );
  INVX1 U643 ( .A(dbg_08[1]), .Y(n664) );
  INVX1 U644 ( .A(dbg_09[1]), .Y(n665) );
  INVX1 U645 ( .A(c_buf_21__4_), .Y(n559) );
  INVX1 U646 ( .A(c_buf_22__4_), .Y(n560) );
  INVX1 U647 ( .A(c_buf_21__0_), .Y(n674) );
  INVX1 U648 ( .A(c_buf_22__0_), .Y(n675) );
  INVX1 U649 ( .A(c_buf_21__3_), .Y(n585) );
  INVX1 U650 ( .A(c_buf_22__3_), .Y(n586) );
  NAND21X1 U651 ( .B(n340), .A(memaddr[14]), .Y(n324) );
  NAND21X1 U652 ( .B(cs_ft[0]), .A(cs_ft[1]), .Y(n202) );
  INVX1 U653 ( .A(cs_ft[3]), .Y(n200) );
  INVX1 U654 ( .A(mcu_psw), .Y(n414) );
  INVX1 U655 ( .A(cs_ft[2]), .Y(n229) );
  INVX1 U656 ( .A(dbg_0a[5]), .Y(n546) );
  INVX1 U657 ( .A(dbg_0b[5]), .Y(n547) );
  INVX1 U658 ( .A(dbg_0a[6]), .Y(n520) );
  INVX1 U659 ( .A(dbg_0b[6]), .Y(n521) );
  INVX1 U660 ( .A(dbg_0a[4]), .Y(n572) );
  INVX1 U661 ( .A(dbg_0b[4]), .Y(n573) );
  INVX1 U662 ( .A(dbg_0a[0]), .Y(n695) );
  INVX1 U663 ( .A(dbg_0b[0]), .Y(n696) );
  INVX1 U664 ( .A(dbg_0a[3]), .Y(n598) );
  INVX1 U665 ( .A(dbg_0b[3]), .Y(n599) );
  INVX1 U666 ( .A(dbg_0a[2]), .Y(n624) );
  INVX1 U667 ( .A(dbg_0b[2]), .Y(n625) );
  INVX1 U668 ( .A(dbg_0a[1]), .Y(n661) );
  INVX1 U669 ( .A(dbg_0b[1]), .Y(n662) );
  NAND21X1 U670 ( .B(d_psrd), .A(n351), .Y(n391) );
  INVX1 U671 ( .A(wr_buf[7]), .Y(n417) );
  INVX1 U672 ( .A(c_buf_18__7_), .Y(n465) );
  INVX1 U673 ( .A(dbg_0f[7]), .Y(n471) );
  INVX1 U674 ( .A(dbg_0c[7]), .Y(n477) );
  INVX1 U675 ( .A(c_buf_20__7_), .Y(n463) );
  INVX1 U676 ( .A(c_buf_17__7_), .Y(n469) );
  INVX1 U677 ( .A(c_buf_19__7_), .Y(n467) );
  INVX1 U678 ( .A(c_buf_16__7_), .Y(n473) );
  INVX1 U679 ( .A(dbg_0d[7]), .Y(n479) );
  NAND43X1 U680 ( .B(pmem_a[11]), .C(pmem_a[10]), .D(adr_p[13]), .A(n785), .Y(
        n784) );
  NOR21XL U681 ( .B(n273), .A(n272), .Y(n280) );
  NOR43XL U682 ( .B(n737), .C(r_multi), .D(n738), .A(pmem_re), .Y(n272) );
  MUX2BXL U683 ( .D0(adr_p[13]), .D1(n783), .S(adr_p[14]), .Y(n279) );
  OAI22X1 U684 ( .A(adr_p[14]), .B(adr_p[13]), .C(pmem_a[9]), .D(n784), .Y(
        n275) );
  INVX1 U685 ( .A(cs_ft[1]), .Y(n94) );
  INVX1 U686 ( .A(cs_ft[0]), .Y(n92) );
  INVX1 U687 ( .A(c_buf_18__5_), .Y(n536) );
  INVX1 U688 ( .A(dbg_0e[7]), .Y(n475) );
  INVX1 U689 ( .A(c_buf_19__5_), .Y(n537) );
  INVX1 U690 ( .A(c_buf_16__5_), .Y(n540) );
  OR2X1 U691 ( .A(cs_ft[3]), .B(n202), .Y(n276) );
  NAND21X1 U692 ( .B(cs_ft[2]), .A(n200), .Y(n97) );
  NAND21X1 U693 ( .B(cs_ft[1]), .A(cs_ft[0]), .Y(n201) );
  NAND21X1 U694 ( .B(n229), .A(cs_ft[3]), .Y(n90) );
  NAND21X1 U695 ( .B(cs_ft[0]), .A(n91), .Y(n107) );
  INVX1 U696 ( .A(n89), .Y(n91) );
  NAND32X1 U697 ( .B(cs_ft[2]), .C(n200), .A(n94), .Y(n89) );
  INVX1 U698 ( .A(wr_buf[0]), .Y(n416) );
  INVX1 U699 ( .A(wr_buf[5]), .Y(n419) );
  INVX1 U700 ( .A(wr_buf[1]), .Y(n423) );
  INVX1 U701 ( .A(wr_buf[3]), .Y(n421) );
  INVX1 U702 ( .A(wr_buf[6]), .Y(n418) );
  INVX1 U703 ( .A(wr_buf[2]), .Y(n422) );
  INVX1 U704 ( .A(wr_buf[4]), .Y(n420) );
  INVX1 U705 ( .A(dbg_0f[5]), .Y(n539) );
  INVX1 U706 ( .A(dbg_0c[5]), .Y(n542) );
  INVX1 U707 ( .A(c_buf_18__6_), .Y(n510) );
  INVX1 U708 ( .A(dbg_0f[6]), .Y(n513) );
  INVX1 U709 ( .A(dbg_0c[6]), .Y(n516) );
  INVX1 U710 ( .A(c_buf_18__4_), .Y(n562) );
  INVX1 U711 ( .A(dbg_0f[4]), .Y(n565) );
  INVX1 U712 ( .A(dbg_0c[4]), .Y(n568) );
  INVX1 U713 ( .A(c_buf_18__0_), .Y(n681) );
  INVX1 U714 ( .A(dbg_0f[0]), .Y(n686) );
  INVX1 U715 ( .A(dbg_0c[0]), .Y(n691) );
  INVX1 U716 ( .A(c_buf_18__3_), .Y(n588) );
  INVX1 U717 ( .A(dbg_0f[3]), .Y(n591) );
  INVX1 U718 ( .A(dbg_0c[3]), .Y(n594) );
  INVX1 U719 ( .A(c_buf_18__2_), .Y(n614) );
  INVX1 U720 ( .A(dbg_0f[2]), .Y(n617) );
  INVX1 U721 ( .A(dbg_0c[2]), .Y(n620) );
  INVX1 U722 ( .A(c_buf_18__1_), .Y(n640) );
  INVX1 U723 ( .A(dbg_0f[1]), .Y(n654) );
  INVX1 U724 ( .A(dbg_0c[1]), .Y(n657) );
  INVX1 U725 ( .A(c_buf_20__5_), .Y(n535) );
  INVX1 U726 ( .A(c_buf_17__5_), .Y(n538) );
  INVX1 U727 ( .A(dbg_0e[5]), .Y(n541) );
  INVX1 U728 ( .A(c_buf_20__6_), .Y(n509) );
  INVX1 U729 ( .A(c_buf_17__6_), .Y(n512) );
  INVX1 U730 ( .A(dbg_0e[6]), .Y(n515) );
  INVX1 U731 ( .A(c_buf_20__4_), .Y(n561) );
  INVX1 U732 ( .A(c_buf_17__4_), .Y(n564) );
  INVX1 U733 ( .A(dbg_0e[4]), .Y(n567) );
  INVX1 U734 ( .A(c_buf_20__0_), .Y(n680) );
  INVX1 U735 ( .A(c_buf_17__0_), .Y(n685) );
  INVX1 U736 ( .A(dbg_0e[0]), .Y(n690) );
  INVX1 U737 ( .A(c_buf_20__3_), .Y(n587) );
  INVX1 U738 ( .A(c_buf_17__3_), .Y(n590) );
  INVX1 U739 ( .A(dbg_0e[3]), .Y(n593) );
  INVX1 U740 ( .A(c_buf_20__2_), .Y(n613) );
  INVX1 U741 ( .A(c_buf_17__2_), .Y(n616) );
  INVX1 U742 ( .A(dbg_0e[2]), .Y(n619) );
  INVX1 U743 ( .A(c_buf_20__1_), .Y(n639) );
  INVX1 U744 ( .A(c_buf_17__1_), .Y(n653) );
  INVX1 U745 ( .A(dbg_0e[1]), .Y(n656) );
  INVX1 U746 ( .A(dbg_0d[5]), .Y(n543) );
  INVX1 U747 ( .A(c_buf_19__6_), .Y(n511) );
  INVX1 U748 ( .A(c_buf_16__6_), .Y(n514) );
  INVX1 U749 ( .A(dbg_0d[6]), .Y(n517) );
  INVX1 U750 ( .A(c_buf_19__4_), .Y(n563) );
  INVX1 U751 ( .A(c_buf_16__4_), .Y(n566) );
  INVX1 U752 ( .A(dbg_0d[4]), .Y(n569) );
  INVX1 U753 ( .A(c_buf_19__0_), .Y(n682) );
  INVX1 U754 ( .A(c_buf_16__0_), .Y(n687) );
  INVX1 U755 ( .A(dbg_0d[0]), .Y(n692) );
  INVX1 U756 ( .A(c_buf_19__3_), .Y(n589) );
  INVX1 U757 ( .A(c_buf_16__3_), .Y(n592) );
  INVX1 U758 ( .A(dbg_0d[3]), .Y(n595) );
  INVX1 U759 ( .A(c_buf_19__2_), .Y(n615) );
  INVX1 U760 ( .A(c_buf_16__2_), .Y(n618) );
  INVX1 U761 ( .A(dbg_0d[2]), .Y(n621) );
  INVX1 U762 ( .A(c_buf_19__1_), .Y(n652) );
  INVX1 U763 ( .A(c_buf_16__1_), .Y(n655) );
  INVX1 U764 ( .A(dbg_0d[1]), .Y(n658) );
  INVX1 U765 ( .A(n291), .Y(n760) );
  XNOR3X1 U766 ( .A(c_adr[2]), .B(c_ptr[2]), .C(n157), .Y(n61) );
  INVX1 U767 ( .A(n158), .Y(n142) );
  NAND21X1 U768 ( .B(n356), .A(c_adr[0]), .Y(n158) );
  XNOR3X1 U769 ( .A(c_adr[4]), .B(c_ptr[4]), .C(n155), .Y(n62) );
  XNOR3X1 U770 ( .A(c_adr[3]), .B(c_ptr[3]), .C(n156), .Y(n63) );
  INVX1 U771 ( .A(c_ptr[0]), .Y(n356) );
  XNOR2XL U772 ( .A(n166), .B(c_adr[5]), .Y(n64) );
  XOR2X1 U773 ( .A(n167), .B(c_adr[6]), .Y(n168) );
  NAND2X1 U774 ( .A(n166), .B(c_adr[5]), .Y(n167) );
  XOR2X1 U775 ( .A(n154), .B(c_adr[7]), .Y(n174) );
  XOR3X1 U776 ( .A(c_adr[1]), .B(c_ptr[1]), .C(n158), .Y(n159) );
  NAND31X1 U777 ( .C(n143), .A(c_adr[5]), .B(n166), .Y(n154) );
  XOR2X1 U778 ( .A(n153), .B(c_adr[8]), .Y(n175) );
  NAND21X1 U779 ( .B(n152), .A(n151), .Y(n153) );
  XOR2X1 U780 ( .A(n150), .B(c_adr[9]), .Y(n178) );
  XOR2X1 U781 ( .A(n356), .B(c_adr[0]), .Y(n209) );
  NAND32X1 U782 ( .B(n145), .C(n180), .A(n179), .Y(n149) );
  INVX1 U783 ( .A(c_adr[10]), .Y(n145) );
  XOR2X1 U784 ( .A(n181), .B(c_adr[10]), .Y(n184) );
  NAND21X1 U785 ( .B(n180), .A(n179), .Y(n181) );
  XOR2X1 U786 ( .A(n149), .B(c_adr[11]), .Y(n187) );
  XOR2X1 U787 ( .A(n148), .B(c_adr[13]), .Y(n195) );
  NAND21X1 U788 ( .B(n148), .A(c_adr[13]), .Y(n147) );
  XOR2X1 U789 ( .A(n190), .B(c_adr[12]), .Y(n192) );
  NAND21X1 U790 ( .B(n189), .A(n188), .Y(n190) );
  INVX1 U791 ( .A(c_adr[2]), .Y(n119) );
  INVX1 U792 ( .A(c_adr[7]), .Y(n152) );
  INVX1 U793 ( .A(c_adr[6]), .Y(n143) );
  INVX1 U794 ( .A(c_adr[9]), .Y(n180) );
  INVX1 U795 ( .A(c_adr[8]), .Y(n144) );
  INVX1 U796 ( .A(c_adr[11]), .Y(n189) );
  INVX1 U797 ( .A(c_adr[12]), .Y(n146) );
  INVX1 U798 ( .A(d_psrd), .Y(n415) );
  INVX1 U799 ( .A(c_adr[13]), .Y(n113) );
  NAND43X1 U800 ( .B(c_ptr[2]), .C(n230), .D(n251), .A(c_ptr[4]), .Y(n238) );
  NAND21X1 U801 ( .B(c_ptr[1]), .A(n356), .Y(n230) );
  INVX1 U802 ( .A(c_ptr[2]), .Y(n373) );
  INVX1 U803 ( .A(c_ptr[3]), .Y(n251) );
  INVX1 U804 ( .A(c_ptr[4]), .Y(n372) );
  NAND21X1 U805 ( .B(n103), .A(n96), .Y(n291) );
  MUX2X1 U806 ( .D0(pmem_q0[7]), .D1(pmem_q1[7]), .S(n105), .Y(n96) );
  NAND21X1 U807 ( .B(n103), .A(n102), .Y(n773) );
  MUX2X1 U808 ( .D0(pmem_q0[1]), .D1(pmem_q1[1]), .S(n105), .Y(n102) );
  NAND21X1 U809 ( .B(n103), .A(n101), .Y(n771) );
  MUX2X1 U810 ( .D0(pmem_q0[2]), .D1(pmem_q1[2]), .S(n105), .Y(n101) );
  NAND21X1 U811 ( .B(n103), .A(n100), .Y(n769) );
  MUX2X1 U812 ( .D0(pmem_q0[3]), .D1(pmem_q1[3]), .S(n105), .Y(n100) );
  NAND21X1 U813 ( .B(n103), .A(n99), .Y(n765) );
  MUX2X1 U814 ( .D0(pmem_q0[5]), .D1(pmem_q1[5]), .S(n105), .Y(n99) );
  NAND21X1 U815 ( .B(n103), .A(n98), .Y(n763) );
  MUX2X1 U816 ( .D0(pmem_q0[6]), .D1(pmem_q1[6]), .S(n105), .Y(n98) );
  OAI22X1 U817 ( .A(pmem_q0[0]), .B(n105), .C(pmem_q1[0]), .D(n104), .Y(n775)
         );
  OAI22X1 U818 ( .A(pmem_q0[4]), .B(n105), .C(pmem_q1[4]), .D(n104), .Y(n767)
         );
  NAND21X1 U819 ( .B(mcu_psw), .A(n360), .Y(n751) );
  INVX1 U820 ( .A(memaddr[13]), .Y(n329) );
  NAND21X1 U821 ( .B(n356), .A(c_ptr[1]), .Y(n375) );
  INVX1 U822 ( .A(n244), .Y(n261) );
  NAND21X1 U823 ( .B(c_ptr[0]), .A(c_ptr[1]), .Y(n244) );
  INVX1 U824 ( .A(n243), .Y(n259) );
  NAND21X1 U825 ( .B(c_ptr[1]), .A(c_ptr[0]), .Y(n243) );
  INVXL U826 ( .A(n281), .Y(n283) );
  AO21XL U827 ( .B(n395), .C(n262), .A(n281), .Y(n311) );
  OAI31XL U828 ( .A(n307), .B(pmem_csb), .C(n281), .D(n108), .Y(n643) );
  NAND21X1 U829 ( .B(pwrdn_rst), .A(n88), .Y(n65) );
  INVXL U830 ( .A(n87), .Y(n85) );
  INVXL U831 ( .A(n382), .Y(n86) );
  OA22XL U832 ( .A(memaddr_c[3]), .B(n63), .C(memaddr_c[2]), .D(n61), .Y(n163)
         );
  INVXL U833 ( .A(memaddr_c[3]), .Y(n410) );
  OAI32XL U834 ( .A(memaddr_c[2]), .B(n119), .C(n118), .D(memaddr_c[3]), .E(
        n431), .Y(n122) );
  MAJ3X1 U835 ( .A(c_adr[1]), .B(c_ptr[1]), .C(n142), .Y(n157) );
  MAJ3X1 U836 ( .A(c_adr[2]), .B(c_ptr[2]), .C(n157), .Y(n156) );
  MAJ3X1 U837 ( .A(c_adr[3]), .B(c_ptr[3]), .C(n156), .Y(n155) );
  MAJ3X1 U838 ( .A(c_adr[4]), .B(c_ptr[4]), .C(n155), .Y(n166) );
  AND2X1 U839 ( .A(c_adr[14]), .B(add_1_root_add_113_2_carry[14]), .Y(N232) );
  XOR2X1 U840 ( .A(add_1_root_add_113_2_carry[14]), .B(c_adr[14]), .Y(N231) );
  AND2X1 U841 ( .A(c_adr[13]), .B(add_1_root_add_113_2_carry[13]), .Y(
        add_1_root_add_113_2_carry[14]) );
  XOR2X1 U842 ( .A(add_1_root_add_113_2_carry[13]), .B(c_adr[13]), .Y(N230) );
  AND2X1 U843 ( .A(c_adr[12]), .B(add_1_root_add_113_2_carry[12]), .Y(
        add_1_root_add_113_2_carry[13]) );
  XOR2X1 U844 ( .A(add_1_root_add_113_2_carry[12]), .B(c_adr[12]), .Y(N229) );
  AND2X1 U845 ( .A(c_adr[11]), .B(add_1_root_add_113_2_carry[11]), .Y(
        add_1_root_add_113_2_carry[12]) );
  XOR2X1 U846 ( .A(add_1_root_add_113_2_carry[11]), .B(c_adr[11]), .Y(N228) );
  AND2X1 U847 ( .A(c_adr[10]), .B(add_1_root_add_113_2_carry[10]), .Y(
        add_1_root_add_113_2_carry[11]) );
  XOR2X1 U848 ( .A(add_1_root_add_113_2_carry[10]), .B(c_adr[10]), .Y(N227) );
  AND2X1 U849 ( .A(c_adr[9]), .B(add_1_root_add_113_2_carry[9]), .Y(
        add_1_root_add_113_2_carry[10]) );
  XOR2X1 U850 ( .A(add_1_root_add_113_2_carry[9]), .B(c_adr[9]), .Y(N226) );
  AND2X1 U851 ( .A(c_adr[8]), .B(add_1_root_add_113_2_carry[8]), .Y(
        add_1_root_add_113_2_carry[9]) );
  XOR2X1 U852 ( .A(add_1_root_add_113_2_carry[8]), .B(c_adr[8]), .Y(N225) );
  AND2X1 U853 ( .A(c_adr[7]), .B(add_1_root_add_113_2_carry[7]), .Y(
        add_1_root_add_113_2_carry[8]) );
  XOR2X1 U854 ( .A(add_1_root_add_113_2_carry[7]), .B(c_adr[7]), .Y(N224) );
  AND2X1 U855 ( .A(c_adr[6]), .B(add_1_root_add_113_2_carry[6]), .Y(
        add_1_root_add_113_2_carry[7]) );
  XOR2X1 U856 ( .A(add_1_root_add_113_2_carry[6]), .B(c_adr[6]), .Y(N223) );
  AND2X1 U857 ( .A(c_adr[5]), .B(add_1_root_add_113_2_carry[5]), .Y(
        add_1_root_add_113_2_carry[6]) );
  XOR2X1 U858 ( .A(add_1_root_add_113_2_carry[5]), .B(c_adr[5]), .Y(N222) );
  OR2X1 U859 ( .A(c_adr[0]), .B(c_ptr[0]), .Y(add_1_root_add_113_2_carry[1])
         );
  XNOR2XL U860 ( .A(c_adr[0]), .B(c_ptr[0]), .Y(N217) );
  OR2X1 U861 ( .A(memaddr[0]), .B(n433), .Y(sub_313_carry[1]) );
  XNOR2XL U862 ( .A(memaddr[0]), .B(n433), .Y(popptr[0]) );
  INVX1 U863 ( .A(wspp_cnt[0]), .Y(N353) );
  OR2X1 U864 ( .A(wspp_cnt[1]), .B(wspp_cnt[0]), .Y(n425) );
  OAI21BBX1 U865 ( .A(wspp_cnt[0]), .B(wspp_cnt[1]), .C(n425), .Y(N354) );
  OR2X1 U866 ( .A(n425), .B(wspp_cnt[2]), .Y(n426) );
  OAI21BBX1 U867 ( .A(n425), .B(wspp_cnt[2]), .C(n426), .Y(N355) );
  OR2X1 U868 ( .A(n426), .B(wspp_cnt[3]), .Y(n427) );
  OAI21BBX1 U869 ( .A(n426), .B(wspp_cnt[3]), .C(n427), .Y(N356) );
  OR2X1 U870 ( .A(n427), .B(wspp_cnt[4]), .Y(n428) );
  OAI21BBX1 U871 ( .A(n427), .B(wspp_cnt[4]), .C(n428), .Y(N357) );
  XNOR2XL U872 ( .A(n428), .B(wspp_cnt[5]), .Y(N358) );
  OR2X1 U873 ( .A(wspp_cnt[5]), .B(n428), .Y(n429) );
  XNOR2XL U874 ( .A(wspp_cnt[6]), .B(n429), .Y(N359) );
  XOR2X1 U875 ( .A(add_255_carry[4]), .B(c_ptr[4]), .Y(N452) );
  OR2X1 U876 ( .A(c_adr[5]), .B(n408), .Y(n436) );
  NAND21X1 U877 ( .B(c_adr[7]), .A(memaddr_c[7]), .Y(n434) );
  NAND21X1 U878 ( .B(c_adr[3]), .A(memaddr_c[3]), .Y(n435) );
  NAND2X1 U879 ( .A(n439), .B(n440), .Y(o_set_hold) );
  NAND4X1 U880 ( .A(n441), .B(n442), .C(n443), .D(n444), .Y(n440) );
  NOR4XL U881 ( .A(n445), .B(memaddr[4]), .C(memaddr[6]), .D(memaddr[5]), .Y(
        n444) );
  OR3XL U882 ( .A(memaddr[8]), .B(memaddr[9]), .C(memaddr[7]), .Y(n445) );
  NOR4XL U883 ( .A(n446), .B(memaddr[12]), .C(memaddr[14]), .D(memaddr[13]), 
        .Y(n443) );
  OR3XL U884 ( .A(memaddr[2]), .B(memaddr[3]), .C(memaddr[1]), .Y(n446) );
  NOR4XL U885 ( .A(n447), .B(memaddr[0]), .C(memaddr[11]), .D(memaddr[10]), 
        .Y(n442) );
  NAND3X1 U886 ( .A(o_inst[6]), .B(o_inst[7]), .C(o_inst[5]), .Y(n447) );
  NOR43XL U887 ( .B(o_inst[0]), .C(o_inst[1]), .D(r_rdy), .A(n448), .Y(n441)
         );
  NAND3X1 U888 ( .A(o_inst[3]), .B(o_inst[4]), .C(o_inst[2]), .Y(n448) );
  NAND4X1 U889 ( .A(n449), .B(n450), .C(n451), .D(n452), .Y(o_inst[7]) );
  NOR4XL U890 ( .A(n453), .B(n454), .C(n455), .D(n456), .Y(n452) );
  OAI222XL U891 ( .A(n457), .B(n417), .C(n458), .D(n459), .E(n460), .F(n461), 
        .Y(n456) );
  OAI222XL U892 ( .A(n462), .B(n463), .C(n464), .D(n465), .E(n466), .F(n467), 
        .Y(n455) );
  OAI222XL U893 ( .A(n468), .B(n469), .C(n470), .D(n471), .E(n472), .F(n473), 
        .Y(n454) );
  OAI222XL U894 ( .A(n474), .B(n475), .C(n476), .D(n477), .E(n478), .F(n479), 
        .Y(n453) );
  AOI211X1 U895 ( .C(dbg_06[7]), .D(n480), .A(n481), .B(n482), .Y(n451) );
  OAI22X1 U896 ( .A(n483), .B(n484), .C(n485), .D(n486), .Y(n482) );
  OAI222XL U897 ( .A(n487), .B(n488), .C(n489), .D(n490), .E(n491), .F(n492), 
        .Y(n481) );
  AOI222XL U898 ( .A(dbg_03[7]), .B(n493), .C(dbg_04[7]), .D(n494), .E(
        dbg_05[7]), .F(n495), .Y(n450) );
  AOI222XL U899 ( .A(rd_buf[7]), .B(n496), .C(dbg_01[7]), .D(n497), .E(
        dbg_02[7]), .F(n498), .Y(n449) );
  NAND4X1 U900 ( .A(n499), .B(n500), .C(n501), .D(n502), .Y(o_inst[6]) );
  NOR4XL U901 ( .A(n503), .B(n504), .C(n505), .D(n506), .Y(n502) );
  OAI222XL U902 ( .A(n457), .B(n418), .C(n458), .D(n507), .E(n460), .F(n508), 
        .Y(n506) );
  OAI222XL U903 ( .A(n462), .B(n509), .C(n464), .D(n510), .E(n466), .F(n511), 
        .Y(n505) );
  OAI222XL U904 ( .A(n468), .B(n512), .C(n470), .D(n513), .E(n472), .F(n514), 
        .Y(n504) );
  OAI222XL U905 ( .A(n474), .B(n515), .C(n476), .D(n516), .E(n478), .F(n517), 
        .Y(n503) );
  AOI211X1 U906 ( .C(dbg_06[6]), .D(n480), .A(n518), .B(n519), .Y(n501) );
  OAI22X1 U907 ( .A(n483), .B(n520), .C(n485), .D(n521), .Y(n519) );
  OAI222XL U908 ( .A(n487), .B(n522), .C(n489), .D(n523), .E(n491), .F(n524), 
        .Y(n518) );
  AOI222XL U909 ( .A(dbg_03[6]), .B(n493), .C(dbg_04[6]), .D(n494), .E(
        dbg_05[6]), .F(n495), .Y(n500) );
  AOI222XL U910 ( .A(rd_buf[6]), .B(n496), .C(dbg_01[6]), .D(n497), .E(
        dbg_02[6]), .F(n498), .Y(n499) );
  NAND4X1 U911 ( .A(n525), .B(n526), .C(n527), .D(n528), .Y(o_inst[5]) );
  NOR4XL U912 ( .A(n529), .B(n530), .C(n531), .D(n532), .Y(n528) );
  OAI222XL U913 ( .A(n457), .B(n419), .C(n458), .D(n533), .E(n460), .F(n534), 
        .Y(n532) );
  OAI222XL U914 ( .A(n462), .B(n535), .C(n464), .D(n536), .E(n466), .F(n537), 
        .Y(n531) );
  OAI222XL U915 ( .A(n468), .B(n538), .C(n470), .D(n539), .E(n472), .F(n540), 
        .Y(n530) );
  OAI222XL U916 ( .A(n474), .B(n541), .C(n476), .D(n542), .E(n478), .F(n543), 
        .Y(n529) );
  AOI211X1 U917 ( .C(dbg_06[5]), .D(n480), .A(n544), .B(n545), .Y(n527) );
  OAI22X1 U918 ( .A(n483), .B(n546), .C(n485), .D(n547), .Y(n545) );
  OAI222XL U919 ( .A(n487), .B(n548), .C(n489), .D(n549), .E(n491), .F(n550), 
        .Y(n544) );
  AOI222XL U920 ( .A(dbg_03[5]), .B(n493), .C(dbg_04[5]), .D(n494), .E(
        dbg_05[5]), .F(n495), .Y(n526) );
  AOI222XL U921 ( .A(rd_buf[5]), .B(n496), .C(dbg_01[5]), .D(n497), .E(
        dbg_02[5]), .F(n498), .Y(n525) );
  NAND4X1 U922 ( .A(n551), .B(n552), .C(n553), .D(n554), .Y(o_inst[4]) );
  NOR4XL U923 ( .A(n555), .B(n556), .C(n557), .D(n558), .Y(n554) );
  OAI222XL U924 ( .A(n457), .B(n420), .C(n458), .D(n559), .E(n460), .F(n560), 
        .Y(n558) );
  OAI222XL U925 ( .A(n462), .B(n561), .C(n464), .D(n562), .E(n466), .F(n563), 
        .Y(n557) );
  OAI222XL U926 ( .A(n468), .B(n564), .C(n470), .D(n565), .E(n472), .F(n566), 
        .Y(n556) );
  OAI222XL U927 ( .A(n474), .B(n567), .C(n476), .D(n568), .E(n478), .F(n569), 
        .Y(n555) );
  AOI211X1 U928 ( .C(dbg_06[4]), .D(n480), .A(n570), .B(n571), .Y(n553) );
  OAI22X1 U929 ( .A(n483), .B(n572), .C(n485), .D(n573), .Y(n571) );
  OAI222XL U930 ( .A(n487), .B(n574), .C(n489), .D(n575), .E(n491), .F(n576), 
        .Y(n570) );
  AOI222XL U931 ( .A(dbg_03[4]), .B(n493), .C(dbg_04[4]), .D(n494), .E(
        dbg_05[4]), .F(n495), .Y(n552) );
  AOI222XL U932 ( .A(rd_buf[4]), .B(n496), .C(dbg_01[4]), .D(n497), .E(
        dbg_02[4]), .F(n498), .Y(n551) );
  NAND4X1 U933 ( .A(n577), .B(n578), .C(n579), .D(n580), .Y(o_inst[3]) );
  NOR4XL U934 ( .A(n581), .B(n582), .C(n583), .D(n584), .Y(n580) );
  OAI222XL U935 ( .A(n457), .B(n421), .C(n458), .D(n585), .E(n460), .F(n586), 
        .Y(n584) );
  OAI222XL U936 ( .A(n462), .B(n587), .C(n464), .D(n588), .E(n466), .F(n589), 
        .Y(n583) );
  OAI222XL U937 ( .A(n468), .B(n590), .C(n470), .D(n591), .E(n472), .F(n592), 
        .Y(n582) );
  OAI222XL U938 ( .A(n474), .B(n593), .C(n476), .D(n594), .E(n478), .F(n595), 
        .Y(n581) );
  AOI211X1 U939 ( .C(dbg_06[3]), .D(n480), .A(n596), .B(n597), .Y(n579) );
  OAI22X1 U940 ( .A(n483), .B(n598), .C(n485), .D(n599), .Y(n597) );
  OAI222XL U941 ( .A(n487), .B(n600), .C(n489), .D(n601), .E(n491), .F(n602), 
        .Y(n596) );
  AOI222XL U942 ( .A(dbg_03[3]), .B(n493), .C(dbg_04[3]), .D(n494), .E(
        dbg_05[3]), .F(n495), .Y(n578) );
  AOI222XL U943 ( .A(rd_buf[3]), .B(n496), .C(dbg_01[3]), .D(n497), .E(
        dbg_02[3]), .F(n498), .Y(n577) );
  NAND4X1 U944 ( .A(n603), .B(n604), .C(n605), .D(n606), .Y(o_inst[2]) );
  NOR4XL U945 ( .A(n607), .B(n608), .C(n609), .D(n610), .Y(n606) );
  OAI222XL U946 ( .A(n457), .B(n422), .C(n458), .D(n611), .E(n460), .F(n612), 
        .Y(n610) );
  OAI222XL U947 ( .A(n462), .B(n613), .C(n464), .D(n614), .E(n466), .F(n615), 
        .Y(n609) );
  OAI222XL U948 ( .A(n468), .B(n616), .C(n470), .D(n617), .E(n472), .F(n618), 
        .Y(n608) );
  OAI222XL U949 ( .A(n474), .B(n619), .C(n476), .D(n620), .E(n478), .F(n621), 
        .Y(n607) );
  AOI211X1 U950 ( .C(dbg_06[2]), .D(n480), .A(n622), .B(n623), .Y(n605) );
  OAI22X1 U951 ( .A(n483), .B(n624), .C(n485), .D(n625), .Y(n623) );
  OAI222XL U952 ( .A(n487), .B(n626), .C(n489), .D(n627), .E(n491), .F(n628), 
        .Y(n622) );
  AOI222XL U953 ( .A(dbg_03[2]), .B(n493), .C(dbg_04[2]), .D(n494), .E(
        dbg_05[2]), .F(n495), .Y(n604) );
  AOI222XL U954 ( .A(rd_buf[2]), .B(n496), .C(dbg_01[2]), .D(n497), .E(
        dbg_02[2]), .F(n498), .Y(n603) );
  NAND4X1 U955 ( .A(n629), .B(n630), .C(n631), .D(n632), .Y(o_inst[1]) );
  NOR4XL U956 ( .A(n633), .B(n634), .C(n635), .D(n636), .Y(n632) );
  OAI222XL U957 ( .A(n457), .B(n423), .C(n458), .D(n637), .E(n460), .F(n638), 
        .Y(n636) );
  OAI222XL U958 ( .A(n462), .B(n639), .C(n464), .D(n640), .E(n466), .F(n652), 
        .Y(n635) );
  OAI222XL U959 ( .A(n468), .B(n653), .C(n470), .D(n654), .E(n472), .F(n655), 
        .Y(n634) );
  OAI222XL U960 ( .A(n474), .B(n656), .C(n476), .D(n657), .E(n478), .F(n658), 
        .Y(n633) );
  AOI211X1 U961 ( .C(dbg_06[1]), .D(n480), .A(n659), .B(n660), .Y(n631) );
  OAI22X1 U962 ( .A(n483), .B(n661), .C(n485), .D(n662), .Y(n660) );
  OAI222XL U963 ( .A(n487), .B(n663), .C(n489), .D(n664), .E(n491), .F(n665), 
        .Y(n659) );
  AOI222XL U964 ( .A(dbg_03[1]), .B(n493), .C(dbg_04[1]), .D(n494), .E(
        dbg_05[1]), .F(n495), .Y(n630) );
  AOI222XL U965 ( .A(rd_buf[1]), .B(n496), .C(dbg_01[1]), .D(n497), .E(
        dbg_02[1]), .F(n498), .Y(n629) );
  NAND4X1 U966 ( .A(n666), .B(n667), .C(n668), .D(n669), .Y(o_inst[0]) );
  NOR4XL U967 ( .A(n670), .B(n671), .C(n672), .D(n673), .Y(n669) );
  OAI222XL U968 ( .A(n457), .B(n416), .C(n458), .D(n674), .E(n460), .F(n675), 
        .Y(n673) );
  NAND2X1 U969 ( .A(n676), .B(n677), .Y(n460) );
  NAND2X1 U970 ( .A(n676), .B(n678), .Y(n458) );
  NAND2X1 U971 ( .A(n676), .B(n679), .Y(n457) );
  OAI222XL U972 ( .A(n462), .B(n680), .C(n464), .D(n681), .E(n466), .F(n682), 
        .Y(n672) );
  NAND2X1 U973 ( .A(n683), .B(n679), .Y(n466) );
  NAND2X1 U974 ( .A(n683), .B(n677), .Y(n464) );
  NAND2X1 U975 ( .A(n676), .B(n684), .Y(n462) );
  AND2X1 U976 ( .A(popptr[4]), .B(popptr[2]), .Y(n676) );
  OAI222XL U977 ( .A(n468), .B(n685), .C(n470), .D(n686), .E(n472), .F(n687), 
        .Y(n671) );
  NAND2X1 U978 ( .A(n683), .B(n684), .Y(n472) );
  NAND2X1 U979 ( .A(n679), .B(n688), .Y(n470) );
  NAND2X1 U980 ( .A(n683), .B(n678), .Y(n468) );
  AND2X1 U981 ( .A(popptr[4]), .B(n689), .Y(n683) );
  OAI222XL U982 ( .A(n474), .B(n690), .C(n476), .D(n691), .E(n478), .F(n692), 
        .Y(n670) );
  NAND2X1 U983 ( .A(n678), .B(n688), .Y(n478) );
  NAND2X1 U984 ( .A(n684), .B(n688), .Y(n476) );
  NAND2X1 U985 ( .A(n677), .B(n688), .Y(n474) );
  AND2X1 U986 ( .A(popptr[3]), .B(popptr[2]), .Y(n688) );
  AOI211X1 U987 ( .C(dbg_06[0]), .D(n480), .A(n693), .B(n694), .Y(n668) );
  OAI22X1 U988 ( .A(n483), .B(n695), .C(n485), .D(n696), .Y(n694) );
  NAND2X1 U989 ( .A(n697), .B(n679), .Y(n485) );
  NAND2X1 U990 ( .A(n697), .B(n677), .Y(n483) );
  OAI222XL U991 ( .A(n487), .B(n698), .C(n489), .D(n699), .E(n491), .F(n700), 
        .Y(n693) );
  NAND2X1 U992 ( .A(n697), .B(n678), .Y(n491) );
  NAND2X1 U993 ( .A(n697), .B(n684), .Y(n489) );
  AND2X1 U994 ( .A(popptr[3]), .B(n689), .Y(n697) );
  NAND2X1 U995 ( .A(n701), .B(n679), .Y(n487) );
  AND2X1 U996 ( .A(n701), .B(n677), .Y(n480) );
  AOI222XL U997 ( .A(dbg_03[0]), .B(n493), .C(dbg_04[0]), .D(n494), .E(
        dbg_05[0]), .F(n495), .Y(n667) );
  AND2X1 U998 ( .A(n701), .B(n678), .Y(n495) );
  AND2X1 U999 ( .A(n701), .B(n684), .Y(n494) );
  NOR3XL U1000 ( .A(popptr[3]), .B(popptr[4]), .C(n689), .Y(n701) );
  INVX1 U1001 ( .A(popptr[2]), .Y(n689) );
  AND2X1 U1002 ( .A(n702), .B(n679), .Y(n493) );
  AND2X1 U1003 ( .A(popptr[1]), .B(popptr[0]), .Y(n679) );
  AOI222XL U1004 ( .A(rd_buf[0]), .B(n496), .C(dbg_01[0]), .D(n497), .E(
        dbg_02[0]), .F(n498), .Y(n666) );
  AND2X1 U1005 ( .A(n702), .B(n677), .Y(n498) );
  AND2X1 U1006 ( .A(popptr[1]), .B(n703), .Y(n677) );
  AND2X1 U1007 ( .A(n702), .B(n678), .Y(n497) );
  NOR2X1 U1008 ( .A(n703), .B(popptr[1]), .Y(n678) );
  INVX1 U1009 ( .A(popptr[0]), .Y(n703) );
  AND2X1 U1010 ( .A(n702), .B(n684), .Y(n496) );
  NOR2X1 U1011 ( .A(popptr[0]), .B(popptr[1]), .Y(n684) );
  NOR3XL U1012 ( .A(popptr[3]), .B(popptr[4]), .C(popptr[2]), .Y(n702) );
  INVX1 U1013 ( .A(n439), .Y(o_bkp_hold) );
  NAND2X1 U1014 ( .A(n704), .B(n705), .Y(n439) );
  NOR4XL U1015 ( .A(n706), .B(n707), .C(n708), .D(n709), .Y(n705) );
  XOR2X1 U1016 ( .A(bkpt_pc[10]), .B(memaddr[10]), .Y(n709) );
  XOR2X1 U1017 ( .A(bkpt_pc[0]), .B(memaddr[0]), .Y(n708) );
  NAND32X1 U1018 ( .B(un_hold), .C(n710), .A(bkpt_ena), .Y(n707) );
  NAND4X1 U1019 ( .A(n711), .B(n712), .C(n713), .D(n714), .Y(n706) );
  XNOR2XL U1020 ( .A(memaddr[11]), .B(bkpt_pc[11]), .Y(n714) );
  XNOR2XL U1021 ( .A(memaddr[12]), .B(bkpt_pc[12]), .Y(n713) );
  XNOR2XL U1022 ( .A(memaddr[13]), .B(bkpt_pc[13]), .Y(n712) );
  XNOR2XL U1023 ( .A(memaddr[14]), .B(bkpt_pc[14]), .Y(n711) );
  NOR4XL U1024 ( .A(n715), .B(n716), .C(n717), .D(n718), .Y(n704) );
  XOR2X1 U1025 ( .A(bkpt_pc[5]), .B(memaddr[5]), .Y(n718) );
  XOR2X1 U1026 ( .A(bkpt_pc[4]), .B(memaddr[4]), .Y(n717) );
  NAND3X1 U1027 ( .A(n719), .B(n720), .C(n721), .Y(n716) );
  XNOR2XL U1028 ( .A(memaddr[2]), .B(bkpt_pc[2]), .Y(n721) );
  XNOR2XL U1029 ( .A(memaddr[3]), .B(bkpt_pc[3]), .Y(n720) );
  XNOR2XL U1030 ( .A(memaddr[1]), .B(bkpt_pc[1]), .Y(n719) );
  NAND4X1 U1031 ( .A(n722), .B(n723), .C(n724), .D(n725), .Y(n715) );
  XNOR2XL U1032 ( .A(memaddr[6]), .B(bkpt_pc[6]), .Y(n725) );
  XNOR2XL U1033 ( .A(memaddr[7]), .B(bkpt_pc[7]), .Y(n724) );
  XNOR2XL U1034 ( .A(memaddr[8]), .B(bkpt_pc[8]), .Y(n723) );
  XNOR2XL U1035 ( .A(memaddr[9]), .B(bkpt_pc[9]), .Y(n722) );
  MUX2IX1 U1036 ( .D0(n727), .D1(n728), .S(n729), .Y(n651) );
  NAND3X1 U1037 ( .A(n730), .B(n88), .C(dummy[0]), .Y(n727) );
  MUX2IX1 U1038 ( .D0(n731), .D1(n732), .S(n729), .Y(n650) );
  AND4X1 U1039 ( .A(dw_ena), .B(sfr_psw), .C(n730), .D(n88), .Y(n729) );
  NAND2X1 U1040 ( .A(dummy[0]), .B(n733), .Y(n732) );
  NAND3X1 U1041 ( .A(n730), .B(n88), .C(dummy[1]), .Y(n731) );
  INVX1 U1042 ( .A(dw_rst), .Y(n730) );
  NAND21X1 U1043 ( .B(wspp_cnt[4]), .A(n739), .Y(n738) );
  OAI21AX1 U1044 ( .B(wspp_cnt[3]), .C(n740), .A(wspp_cnt[6]), .Y(n739) );
  MUX2IX1 U1045 ( .D0(n741), .D1(n742), .S(wspp_cnt[5]), .Y(n737) );
  AND2X1 U1046 ( .A(n743), .B(wspp_cnt[4]), .Y(n742) );
  OAI21X1 U1047 ( .B(wspp_cnt[6]), .C(n740), .A(n743), .Y(n741) );
  NAND2X1 U1048 ( .A(wspp_cnt[6]), .B(wspp_cnt[3]), .Y(n743) );
  MUX2IX1 U1049 ( .D0(n438), .D1(n710), .S(n414), .Y(mempsack) );
  NAND21X1 U1050 ( .B(rd_buf[7]), .A(d_psrd), .Y(d_inst[7]) );
  NAND21X1 U1051 ( .B(rd_buf[6]), .A(n25), .Y(d_inst[6]) );
  NAND21X1 U1052 ( .B(rd_buf[5]), .A(n25), .Y(d_inst[5]) );
  AND2X1 U1053 ( .A(rd_buf[4]), .B(d_psrd), .Y(d_inst[4]) );
  NAND21X1 U1054 ( .B(rd_buf[3]), .A(n25), .Y(d_inst[3]) );
  NAND21X1 U1055 ( .B(rd_buf[2]), .A(n25), .Y(d_inst[2]) );
  NAND21X1 U1056 ( .B(rd_buf[1]), .A(d_psrd), .Y(d_inst[1]) );
  AND2X1 U1057 ( .A(rd_buf[0]), .B(n25), .Y(d_inst[0]) );
  INVX1 U1058 ( .A(n744), .Y(N974) );
  AOI31X1 U1059 ( .A(un_hold), .B(n88), .C(n710), .D(n801), .Y(n744) );
  NOR2X1 U1060 ( .A(n745), .B(srst), .Y(n801) );
  INVX1 U1061 ( .A(r_rdy), .Y(n710) );
  OAI31XL U1062 ( .A(n751), .B(wr_buf[0]), .C(n424), .D(n736), .Y(n750) );
  NAND2X1 U1063 ( .A(n755), .B(n733), .Y(n728) );
  INVX1 U1064 ( .A(dummy[1]), .Y(n733) );
  INVX1 U1065 ( .A(dummy[0]), .Y(n755) );
  OAI31XL U1066 ( .A(n734), .B(n396), .C(n756), .D(n735), .Y(n752) );
  INVX1 U1067 ( .A(n748), .Y(n756) );
  NAND2X1 U1068 ( .A(n753), .B(n754), .Y(n748) );
  NAND2X1 U1069 ( .A(mcu_psw), .B(hit_ps), .Y(n754) );
  NAND4X1 U1070 ( .A(d_hold[3]), .B(d_hold[2]), .C(n757), .D(d_hold[1]), .Y(
        n753) );
  NOR2X1 U1071 ( .A(n745), .B(n758), .Y(n757) );
  INVX1 U1072 ( .A(r_hold_mcu), .Y(n745) );
  NOR41XL U1073 ( .D(n740), .A(wspp_cnt[0]), .B(wspp_cnt[2]), .C(wspp_cnt[1]), 
        .Y(n746) );
  NOR4XL U1074 ( .A(wspp_cnt[3]), .B(wspp_cnt[4]), .C(wspp_cnt[5]), .D(
        wspp_cnt[6]), .Y(n740) );
  OAI21BBX1 U1075 ( .A(N359), .B(n397), .C(n751), .Y(N801) );
  OAI21BBX1 U1076 ( .A(N358), .B(n397), .C(n751), .Y(N800) );
  OAI21BBX1 U1077 ( .A(N357), .B(n397), .C(n751), .Y(N799) );
  AND2X1 U1078 ( .A(N356), .B(n397), .Y(N798) );
  OAI21BBX1 U1079 ( .A(N355), .B(n397), .C(n751), .Y(N797) );
  OAI21BBX1 U1080 ( .A(N354), .B(n397), .C(n751), .Y(N796) );
  OAI21BBX1 U1081 ( .A(N353), .B(n397), .C(n751), .Y(N795) );
  OAI222XL U1082 ( .A(sfr_wdat[7]), .B(n747), .C(n760), .D(n726), .E(
        memdatao[7]), .F(n761), .Y(N793) );
  OAI221X1 U1083 ( .A(memdatao[6]), .B(n761), .C(n398), .D(n417), .E(n762), 
        .Y(N792) );
  EORX1 U1084 ( .A(n394), .B(n763), .C(sfr_wdat[6]), .D(n747), .Y(n762) );
  OAI221X1 U1085 ( .A(memdatao[5]), .B(n761), .C(n398), .D(n418), .E(n764), 
        .Y(N791) );
  EORX1 U1086 ( .A(n394), .B(n765), .C(sfr_wdat[5]), .D(n747), .Y(n764) );
  OAI221X1 U1087 ( .A(memdatao[4]), .B(n761), .C(n398), .D(n419), .E(n766), 
        .Y(N790) );
  EORX1 U1088 ( .A(n394), .B(n767), .C(sfr_wdat[4]), .D(n747), .Y(n766) );
  OAI221X1 U1089 ( .A(memdatao[3]), .B(n761), .C(n398), .D(n420), .E(n768), 
        .Y(N789) );
  EORX1 U1090 ( .A(n394), .B(n769), .C(sfr_wdat[3]), .D(n747), .Y(n768) );
  OAI221X1 U1091 ( .A(memdatao[2]), .B(n761), .C(n398), .D(n421), .E(n770), 
        .Y(N788) );
  EORX1 U1092 ( .A(n394), .B(n771), .C(sfr_wdat[2]), .D(n747), .Y(n770) );
  OAI221X1 U1093 ( .A(memdatao[1]), .B(n761), .C(n398), .D(n422), .E(n772), 
        .Y(N787) );
  EORX1 U1094 ( .A(n394), .B(n773), .C(sfr_wdat[1]), .D(n747), .Y(n772) );
  OAI221X1 U1095 ( .A(memdatao[0]), .B(n761), .C(n398), .D(n423), .E(n774), 
        .Y(N786) );
  EORX1 U1096 ( .A(n394), .B(n775), .C(sfr_wdat[0]), .D(n747), .Y(n774) );
  NAND2X1 U1097 ( .A(n395), .B(mcu_psw), .Y(n761) );
  NOR2X1 U1098 ( .A(cs_ft[1]), .B(cs_ft[0]), .Y(n759) );
  MUX2IX1 U1099 ( .D0(n776), .D1(n777), .S(pmem_a[8]), .Y(N759) );
  AOI21X1 U1100 ( .B(n778), .C(n779), .A(N757), .Y(n777) );
  NAND3X1 U1101 ( .A(pmem_a[6]), .B(n778), .C(pmem_a[7]), .Y(n776) );
  MUX2BXL U1102 ( .D0(N757), .D1(n780), .S(n779), .Y(N758) );
  INVX1 U1103 ( .A(pmem_a[7]), .Y(n779) );
  NAND2X1 U1104 ( .A(pmem_a[6]), .B(n778), .Y(n780) );
  NOR21XL U1105 ( .B(n778), .A(pmem_a[6]), .Y(N757) );
  NOR2X1 U1106 ( .A(n424), .B(n398), .Y(n778) );
  NAND2X1 U1107 ( .A(n781), .B(n782), .Y(n749) );
  NOR4XL U1108 ( .A(wr_buf[7]), .B(wr_buf[6]), .C(wr_buf[5]), .D(wr_buf[4]), 
        .Y(n782) );
  NOR4XL U1109 ( .A(wr_buf[3]), .B(wr_buf[2]), .C(wr_buf[1]), .D(wr_buf[0]), 
        .Y(n781) );
  NAND21X1 U1110 ( .B(n784), .A(pmem_a[9]), .Y(n783) );
  NOR4XL U1111 ( .A(pmem_a[15]), .B(pmem_a[14]), .C(pmem_a[13]), .D(pmem_a[12]), .Y(n785) );
  XNOR2XL U1112 ( .A(N219), .B(n411), .Y(n788) );
  XNOR2XL U1113 ( .A(N218), .B(n412), .Y(n787) );
  XNOR2XL U1114 ( .A(N217), .B(n413), .Y(n786) );
  XNOR2XL U1115 ( .A(N223), .B(n407), .Y(n792) );
  XNOR2XL U1116 ( .A(N222), .B(n408), .Y(n791) );
  XNOR2XL U1117 ( .A(N221), .B(n409), .Y(n790) );
  XNOR2XL U1118 ( .A(N220), .B(n410), .Y(n789) );
  XNOR2XL U1119 ( .A(N227), .B(n403), .Y(n796) );
  XNOR2XL U1120 ( .A(N226), .B(n404), .Y(n795) );
  XNOR2XL U1121 ( .A(N225), .B(n405), .Y(n794) );
  XNOR2XL U1122 ( .A(N224), .B(n406), .Y(n793) );
  XNOR2XL U1123 ( .A(N231), .B(n399), .Y(n800) );
  XNOR2XL U1124 ( .A(N230), .B(n400), .Y(n799) );
  XNOR2XL U1125 ( .A(N229), .B(n401), .Y(n798) );
  XNOR2XL U1126 ( .A(N228), .B(n402), .Y(n797) );
  AND2X1 U1127 ( .A(d_hold[2]), .B(n88), .Y(N154) );
  AND2X1 U1128 ( .A(d_hold[1]), .B(n88), .Y(N153) );
  NOR2X1 U1129 ( .A(srst), .B(n758), .Y(N152) );
  INVX1 U1130 ( .A(d_hold[0]), .Y(n758) );
  INVX1 U1131 ( .A(n438), .Y(o_ofs_inc) );
endmodule


module ictlr_a0_DW01_inc_2 ( A, SUM );
  input [14:0] A;
  output [14:0] SUM;

  wire   [14:2] carry;

  HAD1X1 U1_1_13 ( .A(A[13]), .B(carry[13]), .CO(carry[14]), .SO(SUM[13]) );
  HAD1X1 U1_1_12 ( .A(A[12]), .B(carry[12]), .CO(carry[13]), .SO(SUM[12]) );
  HAD1X1 U1_1_11 ( .A(A[11]), .B(carry[11]), .CO(carry[12]), .SO(SUM[11]) );
  HAD1X1 U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .SO(SUM[10]) );
  HAD1X1 U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .SO(SUM[9]) );
  HAD1X1 U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .SO(SUM[8]) );
  HAD1X1 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .SO(SUM[7]) );
  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  XOR2X1 U1 ( .A(carry[14]), .B(A[14]), .Y(SUM[14]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module ictlr_a0_DW01_inc_1 ( A, SUM );
  input [14:0] A;
  output [14:0] SUM;

  wire   [14:2] carry;

  HAD1X1 U1_1_13 ( .A(A[13]), .B(carry[13]), .CO(carry[14]), .SO(SUM[13]) );
  HAD1X1 U1_1_12 ( .A(A[12]), .B(carry[12]), .CO(carry[13]), .SO(SUM[12]) );
  HAD1X1 U1_1_11 ( .A(A[11]), .B(carry[11]), .CO(carry[12]), .SO(SUM[11]) );
  HAD1X1 U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .SO(SUM[10]) );
  HAD1X1 U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .SO(SUM[9]) );
  HAD1X1 U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .SO(SUM[8]) );
  HAD1X1 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .SO(SUM[7]) );
  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  XOR2X1 U1 ( .A(carry[14]), .B(A[14]), .Y(SUM[14]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_3 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_4 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_5 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_6 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_7 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_8 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_9 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_10 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_11 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_12 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_13 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_14 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_15 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_16 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_17 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_18 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_19 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_20 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_21 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_22 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_23 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_24 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_25 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_26 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_27 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_28 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_29 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ictlr_a0_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module mcu51_a0 ( bclki2c, pc_ini, slp2wakeup, r_hold_mcu, wdt_slow, wdtov, 
        mdubsy, cs_run, t0_intr, clki2c, clkmdu, clkur0, clktm0, clktm1, 
        clkwdt, i2c_autoack, i2c_con_ens1, clkcpu, clkper, reset, ro, port0i, 
        exint_9, exint, clkcpuen, clkperen, port0o, port0ff, rxd0o, txd0, 
        rxd0i, rxd0oe, scli, sdai, sclo, sdao, waitstaten, mempsack, memack, 
        memdatai, memdatao, memaddr, mempswr, mempsrd, memwr, memrd, 
        memdatao_comb, memaddr_comb, mempswr_comb, mempsrd_comb, memwr_comb, 
        memrd_comb, ramdatai, ramdatao, ramaddr, ramwe, ramoe, dbgpo, sfrack, 
        sfrdatai, sfrdatao, sfraddr, sfrwe, sfroe, esfrm_wrdata, esfrm_addr, 
        esfrm_we, esfrm_oe, esfrm_rddata );
  input [15:0] pc_ini;
  output [1:0] wdtov;
  input [7:0] port0i;
  input [7:0] exint;
  output [7:0] port0o;
  output [7:0] port0ff;
  input [7:0] memdatai;
  output [7:0] memdatao;
  output [15:0] memaddr;
  output [7:0] memdatao_comb;
  output [15:0] memaddr_comb;
  input [7:0] ramdatai;
  output [7:0] ramdatao;
  output [7:0] ramaddr;
  output [31:0] dbgpo;
  input [7:0] sfrdatai;
  output [7:0] sfrdatao;
  output [6:0] sfraddr;
  input [7:0] esfrm_wrdata;
  input [6:0] esfrm_addr;
  output [7:0] esfrm_rddata;
  input bclki2c, slp2wakeup, r_hold_mcu, wdt_slow, clki2c, clkmdu, clkur0,
         clktm0, clktm1, clkwdt, i2c_autoack, clkcpu, clkper, reset, exint_9,
         rxd0i, scli, sdai, mempsack, memack, sfrack, esfrm_we, esfrm_oe;
  output mdubsy, cs_run, t0_intr, i2c_con_ens1, ro, clkcpuen, clkperen, rxd0o,
         txd0, rxd0oe, sclo, sdao, waitstaten, mempswr, mempsrd, memwr, memrd,
         mempswr_comb, mempsrd_comb, memwr_comb, memrd_comb, ramwe, ramoe,
         sfrwe, sfroe;
  wire   n102, n103, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18,
         N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32,
         N33, N34, t0_tf1, t1_tf1, t0_tr1, t1_tr1, stop_flag, idle_flag,
         isfrwait, sfroe_s, sfroe_mcu51_per, sfrwe_s, sfrwe_mcu51_per,
         newinstr, intcall_int, cpu_resume, rmwinstr, pmw, p2sel, gf0, c, ac,
         ov, f0, f1, p, rsttowdt, rsttosrst, rst, int0ff, int1ff, rxd0ff,
         sdaiff, rsttowdtff, rsttosrstff, resetff, smod, ip0wdts, wdt_tm, bd,
         ie0, it0, ie1, it1, iex2, iex3, iex4, iex5, iex6, iex7, iex8, iex9,
         isr_tm, i2c_int, i2ccon_o_7, tf1_gate, riti0_gate, iex7_gate,
         iex2_gate, srstflag, int_vect_8b, int_vect_93, int_vect_9b,
         int_vect_a3, wdts, srst, pmuintreq_rev, pmuintreq, t1ov, t0ack, t1ack,
         isr_irq, int0ack, int1ack, iex7ack, iex2ack, iex3ack, iex4ack,
         iex5ack, iex6ack, iex8ack, iex9ack, n6, n7, n8, n9, n10, n11, n1, n2,
         n3, n4, n5, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n28, n38, n40, n41, n42, n43, n44, n46, n48, n50,
         n51, n53, n54, n55, n56, n58, n60, n62, n64, n66, n68, n70, n72, n74,
         n75, n76, n77, n78, n79, n81, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2,
         SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4,
         SYNOPSYS_UNCONNECTED_5;
  wire   [13:0] timer_1ms;
  wire   [5:0] ien2;
  wire   [6:0] ramsfraddr;
  wire   [4:0] intvect_int;
  wire   [7:0] ckcon;
  wire   [7:0] dph;
  wire   [7:0] dpl;
  wire   [3:0] dps;
  wire   [7:0] p2;
  wire   [5:0] dpc;
  wire   [7:0] sp;
  wire   [7:0] acc_s;
  wire   [7:0] b;
  wire   [1:0] rs;
  wire   [7:0] arcon;
  wire   [7:0] md0;
  wire   [7:0] md1;
  wire   [7:0] md2;
  wire   [7:0] md3;
  wire   [7:0] md4;
  wire   [7:0] md5;
  wire   [3:0] t0_tmod;
  wire   [7:0] tl0;
  wire   [7:0] th0;
  wire   [3:0] t1_tmod;
  wire   [7:0] tl1;
  wire   [7:0] th1;
  wire   [7:0] wdtrel;
  wire   [6:5] t2con;
  wire   [7:0] s0con;
  wire   [7:0] s0buf;
  wire   [7:0] s0rell;
  wire   [7:0] s0relh;
  wire   [7:0] ien0;
  wire   [5:0] ien1;
  wire   [5:0] ip0;
  wire   [5:0] ip1;
  wire   [7:0] i2cdat_o;
  wire   [7:0] i2cadr_o;
  wire   [5:0] i2ccon_o;
  wire   [7:0] i2csta_o;
  wire   [3:0] isreg;

  mcu51_cpu_a0 u_cpu ( .clkcpu(clkcpu), .rst(dbgpo[22]), .mempsack(mempsack), 
        .memack(memack), .memdatai(memdatai), .memaddr(memaddr), .mempsrd(
        mempsrd), .mempswr(mempswr), .memrd(memrd), .memwr(memwr), 
        .memaddr_comb(memaddr_comb), .mempsrd_comb(mempsrd_comb), 
        .mempswr_comb(mempswr_comb), .memrd_comb(memrd_comb), .memwr_comb(
        memwr_comb), .cpu_hold(r_hold_mcu), .cpu_resume(cpu_resume), .irq(
        dbgpo[20]), .intvect(intvect_int), .intcall(intcall_int), .retiinstr(
        dbgpo[21]), .newinstr(newinstr), .rmwinstr(rmwinstr), .waitstaten(
        waitstaten), .ramdatai(ramdatai), .sfrdatai(esfrm_rddata), 
        .ramsfraddr({SYNOPSYS_UNCONNECTED_1, ramsfraddr}), .ramdatao(memdatao), 
        .ramoe(), .ramwe(), .sfroe(sfroe_s), .sfrwe(sfrwe_s), .sfroe_r(), 
        .sfrwe_r(), .sfroe_comb_s(), .sfrwe_comb_s(), .pc_o(dbgpo[15:0]), 
        .pc_ini(pc_ini), .cs_run(cs_run), .instr(dbgpo[31:24]), .codefetch_s(), 
        .sfrack(sfrack), .ramsfraddr_comb(ramaddr), .ramdatao_comb(ramdatao), 
        .ramoe_comb(ramoe), .ramwe_comb(ramwe), .ckcon(ckcon), .pmw(pmw), 
        .p2sel(p2sel), .gf0(gf0), .stop(stop_flag), .idle(idle_flag), .acc(
        acc_s), .b(b), .rs(rs), .c(c), .ac(ac), .ov(ov), .p(p), .f0(f0), .f1(
        f1), .dph(dph), .dpl(dpl), .dps(dps), .dpc(dpc), .p2(p2), .sp(sp) );
  syncneg_a0 u_syncneg ( .clk(clkper), .reset(n75), .rsttowdt(rsttowdt), 
        .rsttosrst(rsttosrst), .rst(rst), .int0(exint[0]), .int1(exint[1]), 
        .port0i(port0i), .rxd0i(rxd0i), .sdai(sdai), .int0ff(int0ff), .int1ff(
        int1ff), .port0ff(port0ff), .t0ff(), .t1ff(), .rxd0ff(rxd0ff), 
        .sdaiff(sdaiff), .rsttowdtff(rsttowdtff), .rsttosrstff(rsttosrstff), 
        .rstff(n102), .resetff(resetff) );
  sfrmux_a0 u_sfrmux ( .isfrwait(isfrwait), .sfraddr({n56, n103, n53, n50, n38, 
        n43, sfraddr[0]}), .c(c), .ac(ac), .f0(f0), .rs(rs), .ov(ov), .f1(f1), 
        .p(p), .acc(acc_s), .b(b), .dpl(dpl), .dph(dph), .dps(dps), .dpc(dpc), 
        .p2(p2), .sp(sp), .smod(smod), .pmw(pmw), .p2sel(p2sel), .gf0(gf0), 
        .stop(stop_flag), .idle(idle_flag), .ckcon(ckcon), .port0(port0o), 
        .port0ff(port0ff), .rmwinstr(rmwinstr), .arcon(arcon), .md0(md0), 
        .md1(md1), .md2(md2), .md3(md3), .md4(md4), .md5(md5), .t0_tmod(
        t0_tmod), .t0_tf0(dbgpo[17]), .t0_tf1(t0_tf1), .t0_tr0(dbgpo[16]), 
        .t0_tr1(t0_tr1), .tl0(tl0), .th0(th0), .t1_tmod(t1_tmod), .t1_tf1(
        t1_tf1), .t1_tr1(t1_tr1), .tl1(tl1), .th1(th1), .wdtrel(wdtrel), 
        .ip0wdts(ip0wdts), .wdt_tm(wdt_tm), .t2con({1'b0, t2con, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .s0con(s0con), .s0buf(s0buf), .s0rell(s0rell), 
        .s0relh(s0relh), .bd(bd), .ie0(ie0), .it0(it0), .ie1(ie1), .it1(it1), 
        .iex2(iex2), .iex3(iex3), .iex4(iex4), .iex5(iex5), .iex6(iex6), 
        .iex7(iex7), .iex8(iex8), .iex9(iex9), .iex10(1'b0), .iex11(1'b0), 
        .iex12(1'b0), .ien0({ien0[7], 1'b0, ien0[5:0]}), .ien1(ien1), .ien2(
        ien2), .ip0(ip0), .ip1(ip1), .isr_tm(isr_tm), .i2c_int(i2c_int), 
        .i2cdat_o(i2cdat_o), .i2cadr_o(i2cadr_o), .i2ccon_o({i2ccon_o_7, 
        i2c_con_ens1, i2ccon_o}), .i2csta_o({i2csta_o[7:3], 1'b0, 1'b0, 1'b0}), 
        .sfrdatai(sfrdatai), .tf1_gate(tf1_gate), .riti0_gate(riti0_gate), 
        .iex7_gate(iex7_gate), .iex2_gate(iex2_gate), .srstflag(srstflag), 
        .int_vect_8b(int_vect_8b), .int_vect_93(int_vect_93), .int_vect_9b(
        int_vect_9b), .int_vect_a3(int_vect_a3), .ext_sfr_sel(), .sfrdatao(
        esfrm_rddata) );
  pmurstctrl_a0 u_pmurstctrl ( .resetff(resetff), .wdts(wdts), .srst(srst), 
        .pmuintreq(pmuintreq_rev), .stop(stop_flag), .idle(idle_flag), 
        .clkcpu_en(clkcpuen), .clkper_en(clkperen), .cpu_resume(cpu_resume), 
        .rsttowdt(rsttowdt), .rsttosrst(rsttosrst), .rst(rst) );
  wakeupctrl_a0 u_wakeupctrl ( .irq(dbgpo[20]), .int0ff(exint[0]), .int1ff(
        exint[1]), .it0(it0), .it1(it1), .isreg(isreg), .intprior0({ip0[2], 
        ip0[0]}), .intprior1({ip1[2], ip1[0]}), .eal(ien0[7]), .eint0(ien0[0]), 
        .eint1(ien0[2]), .pmuintreq(pmuintreq) );
  mdu_a0 u_mdu ( .clkper(clkmdu), .rst(n77), .mdubsy(mdubsy), .sfrdatai({
        sfrdatao[7], n20, sfrdatao[5:0]}), .sfraddr({n58, n5, n53, n51, n46, 
        n44, n41}), .sfrwe(sfrwe_mcu51_per), .sfroe(sfroe_mcu51_per), .arcon(
        arcon), .md0(md0), .md1(md1), .md2(md2), .md3(md3), .md4(md4), .md5(
        md5) );
  ports_a0 u_ports ( .clkper(clkper), .rst(dbgpo[22]), .port0(port0o), 
        .sfrdatai({sfrdatao[7], n20, n25, n22, sfrdatao[3:0]}), .sfraddr({n58, 
        n103, n54, n51, n15, n17, n4}), .sfrwe(n13) );
  serial0_a0 u_serial0 ( .t_shift_clk(), .r_shift_clk(), .clkper(clkur0), 
        .rst(n81), .newinstr(newinstr), .rxd0ff(rxd0ff), .t1ov(t1ov), .rxd0o(
        rxd0o), .rxd0oe(rxd0oe), .txd0(txd0), .sfrdatai({n21, sfrdatao[6:4], 
        n18, n24, n23, n19}), .sfraddr({sfraddr[6], n55, n53, n50, n46, 
        sfraddr[1], n3}), .sfrwe(n13), .s0con(s0con), .s0buf(s0buf), .s0rell(
        s0rell), .s0relh(s0relh), .smod(smod), .bd(bd) );
  timer0_a0 u_timer0 ( .clkper(clktm0), .rst(dbgpo[22]), .newinstr(newinstr), 
        .t0ff(1'b0), .t0ack(t0ack), .t1ack(t1ack), .int0ff(int0ff), .t0_tf0(
        dbgpo[17]), .t0_tf1(t0_tf1), .sfrdatai({n21, sfrdatao[6:4], n18, 
        sfrdatao[2], n23, n19}), .sfraddr({n58, n55, n54, n51, n15, n17, 
        sfraddr[0]}), .sfrwe(n13), .t0_tmod(t0_tmod), .t0_tr0(dbgpo[16]), 
        .t0_tr1(t0_tr1), .tl0(tl0), .th0(th0) );
  timer1_a0 u_timer1 ( .clkper(clktm1), .rst(dbgpo[22]), .newinstr(newinstr), 
        .t1ff(1'b0), .t1ack(t1ack), .int1ff(int1ff), .t1_tf1(t1_tf1), .t1ov(
        t1ov), .sfrdatai({sfrdatao[7:4], n18, sfrdatao[2], n23, n19}), 
        .sfraddr({n58, n5, n54, n51, sfraddr[2], n17, n4}), .sfrwe(n13), 
        .t1_tmod(t1_tmod), .t1_tr1(t1_tr1), .tl1(tl1), .th1(th1) );
  watchdog_a0 u_watchdog ( .wdt_slow(wdt_slow), .clkwdt(clkwdt), .clkper(
        clkper), .resetff(rsttowdtff), .newinstr(newinstr), .wdts_s(wdtov), 
        .wdts(wdts), .ip0wdts(ip0wdts), .wdt_tm(wdt_tm), .sfrdatai({
        sfrdatao[7:6], n25, n22, sfrdatao[3:0]}), .sfraddr({sfraddr[6], n5, 
        n54, sfraddr[3:1], n3}), .sfrwe(n13), .wdtrel(wdtrel) );
  isr_a0 u_isr ( .clkper(clkper), .rst(n78), .intcall(intcall_int), 
        .retiinstr(dbgpo[21]), .int_vect_03(ie0), .int_vect_0b(dbgpo[17]), 
        .t0ff(1'b0), .int_vect_13(ie1), .int_vect_1b(tf1_gate), .t1ff(1'b0), 
        .int_vect_23(riti0_gate), .i2c_int(i2c_int), .rxd0ff(rxd0ff), 
        .int_vect_43(iex7_gate), .sdaiff(sdaiff), .int_vect_4b(iex2_gate), 
        .int_vect_53(iex3), .int_vect_5b(iex4), .int_vect_63(iex5), 
        .int_vect_6b(iex6), .int_vect_8b(int_vect_8b), .int_vect_93(
        int_vect_93), .int_vect_9b(int_vect_9b), .int_vect_a3(int_vect_a3), 
        .int_vect_ab(1'b0), .irq(isr_irq), .intvect(intvect_int), .int_ack_03(
        int0ack), .int_ack_0b(t0ack), .int_ack_13(int1ack), .int_ack_1b(t1ack), 
        .int_ack_43(iex7ack), .int_ack_4b(iex2ack), .int_ack_53(iex3ack), 
        .int_ack_5b(iex4ack), .int_ack_63(iex5ack), .int_ack_6b(iex6ack), 
        .int_ack_8b(iex8ack), .int_ack_93(iex9ack), .int_ack_9b(), 
        .int_ack_a3(), .int_ack_ab(), .is_reg(isreg), .ip0(ip0), .ip1(ip1), 
        .ien0({ien0[7], SYNOPSYS_UNCONNECTED_2, ien0[5:0]}), .ien1(ien1), 
        .ien2(ien2), .isr_tm(isr_tm), .sfraddr({n58, n55, n54, sfraddr[3], n46, 
        n44, n4}), .sfrdatai({sfrdatao[7], n20, n25, sfrdatao[4:0]}), .sfrwe(
        n13) );
  extint_a0 u_extint ( .clkper(clkper), .rst(n79), .newinstr(newinstr), 
        .int0ff(int0ff), .int0ack(int0ack), .int1ff(int1ff), .int1ack(int1ack), 
        .int2ff(exint[2]), .iex2ack(iex2ack), .int3ff(exint[3]), .iex3ack(
        iex3ack), .int4ff(exint[4]), .iex4ack(iex4ack), .int5ff(exint[5]), 
        .iex5ack(iex5ack), .int6ff(exint[6]), .iex6ack(iex6ack), .int7ff(
        exint[7]), .iex7ack(iex7ack), .int8ff(n11), .iex8ack(iex8ack), 
        .int9ff(exint_9), .iex9ack(iex9ack), .ie0(ie0), .it0(it0), .ie1(ie1), 
        .it1(it1), .i2fr(t2con[5]), .iex2(iex2), .i3fr(t2con[6]), .iex3(iex3), 
        .iex4(iex4), .iex5(iex5), .iex6(iex6), .iex7(iex7), .iex8(iex8), 
        .iex9(iex9), .iex10(), .iex11(), .iex12(), .sfraddr({n58, n5, n54, n50, 
        n15, n43, n3}), .sfrdatai({sfrdatao[7], n20, sfrdatao[5], n22, n18, 
        n24, sfrdatao[1], n19}), .sfrwe(n13) );
  i2c_a0 u_i2c ( .clk(clki2c), .rst(n81), .bclksel(bclki2c), .scli(scli), 
        .sdai(sdai), .sclo(sclo), .sdao(sdao), .intack(i2c_autoack), .si(
        i2c_int), .sfrwe(sfrwe_mcu51_per), .sfraddr({sfraddr[6], n55, n54, n51, 
        n15, n44, n41}), .sfrdatai({sfrdatao[7], n20, n25, sfrdatao[4:3], n24, 
        sfrdatao[1:0]}), .i2cdat_o(i2cdat_o), .i2cadr_o(i2cadr_o), .i2ccon_o({
        i2ccon_o_7, i2c_con_ens1, i2ccon_o}), .i2csta_o({i2csta_o[7:3], 
        SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5}) );
  softrstctrl_a0 u_softrstctrl ( .clkcpu(clkcpu), .resetff(rsttosrstff), 
        .newinstr(newinstr), .srstreq(srst), .srstflag(srstflag), .sfrdatai({
        sfrdatao[7], n20, n25, n22, sfrdatao[3:0]}), .sfraddr({n58, n5, n54, 
        n51, sfraddr[2], n43, n41}), .sfrwe(n13) );
  mcu51_a0_DW01_inc_0 add_268 ( .A(timer_1ms), .SUM({N20, N19, N18, N17, N16, 
        N15, N14, N13, N12, N11, N10, N9, N8, N7}) );
  DFFQX1 timer_1ms_reg_13_ ( .D(N34), .C(clkper), .Q(timer_1ms[13]) );
  DFFQX1 timer_1ms_reg_8_ ( .D(N29), .C(clkper), .Q(timer_1ms[8]) );
  DFFQX1 timer_1ms_reg_9_ ( .D(N30), .C(clkper), .Q(timer_1ms[9]) );
  DFFQX1 timer_1ms_reg_10_ ( .D(N31), .C(clkper), .Q(timer_1ms[10]) );
  DFFQX1 timer_1ms_reg_11_ ( .D(N32), .C(clkper), .Q(timer_1ms[11]) );
  DFFQX1 timer_1ms_reg_12_ ( .D(N33), .C(clkper), .Q(timer_1ms[12]) );
  DFFQX1 timer_1ms_reg_5_ ( .D(N26), .C(clkper), .Q(timer_1ms[5]) );
  DFFQX1 timer_1ms_reg_6_ ( .D(N27), .C(clkper), .Q(timer_1ms[6]) );
  DFFQX1 timer_1ms_reg_7_ ( .D(N28), .C(clkper), .Q(timer_1ms[7]) );
  DFFQX1 timer_1ms_reg_4_ ( .D(N25), .C(clkper), .Q(timer_1ms[4]) );
  DFFQX1 timer_1ms_reg_3_ ( .D(N24), .C(clkper), .Q(timer_1ms[3]) );
  DFFQX1 timer_1ms_reg_2_ ( .D(N23), .C(clkper), .Q(timer_1ms[2]) );
  DFFQX1 timer_1ms_reg_1_ ( .D(N22), .C(clkper), .Q(timer_1ms[1]) );
  DFFQX1 timer_1ms_reg_0_ ( .D(N21), .C(clkper), .Q(timer_1ms[0]) );
  MUX2IX1 U3 ( .D0(esfrm_addr[1]), .D1(ramsfraddr[1]), .S(n89), .Y(n26) );
  BUFX3 U4 ( .A(n14), .Y(n1) );
  BUFX3 U5 ( .A(n14), .Y(n2) );
  INVXL U6 ( .A(isfrwait), .Y(n14) );
  MUX2X1 U7 ( .D0(esfrm_addr[0]), .D1(ramsfraddr[0]), .S(n89), .Y(sfraddr[0])
         );
  MUX2IX1 U8 ( .D0(esfrm_addr[6]), .D1(ramsfraddr[6]), .S(n89), .Y(n87) );
  MUX2IX1 U9 ( .D0(esfrm_addr[5]), .D1(ramsfraddr[5]), .S(n89), .Y(n86) );
  INVX1 U10 ( .A(n48), .Y(sfraddr[2]) );
  INVX1 U11 ( .A(n18), .Y(n66) );
  INVXL U12 ( .A(n42), .Y(n3) );
  INVXL U13 ( .A(n42), .Y(n4) );
  INVXL U14 ( .A(n86), .Y(n5) );
  AO21XL U15 ( .B(n92), .C(n76), .A(esfrm_we), .Y(sfrwe) );
  INVX1 U16 ( .A(sfrwe_mcu51_per), .Y(n12) );
  INVX1 U17 ( .A(n12), .Y(n13) );
  INVX3 U18 ( .A(isfrwait), .Y(n89) );
  NAND21X2 U19 ( .B(esfrm_oe), .A(n91), .Y(isfrwait) );
  INVXL U20 ( .A(n48), .Y(n15) );
  INVX1 U21 ( .A(n6), .Y(n40) );
  INVX1 U22 ( .A(n40), .Y(n16) );
  INVXL U23 ( .A(n26), .Y(n17) );
  INVX1 U24 ( .A(n26), .Y(n43) );
  INVX1 U25 ( .A(n28), .Y(n53) );
  INVXL U26 ( .A(n26), .Y(sfraddr[1]) );
  INVX3 U27 ( .A(n85), .Y(n50) );
  INVXL U28 ( .A(n28), .Y(sfraddr[4]) );
  INVXL U29 ( .A(n85), .Y(sfraddr[3]) );
  INVXL U30 ( .A(n28), .Y(n54) );
  INVXL U31 ( .A(n85), .Y(n51) );
  MUX2BXL U32 ( .D0(esfrm_wrdata[3]), .D1(n88), .S(n2), .Y(n18) );
  MUX2XL U33 ( .D0(esfrm_wrdata[0]), .D1(memdatao[0]), .S(n2), .Y(n19) );
  MUX2XL U34 ( .D0(esfrm_wrdata[6]), .D1(memdatao[6]), .S(n2), .Y(n20) );
  MUX2XL U35 ( .D0(esfrm_wrdata[7]), .D1(memdatao[7]), .S(n2), .Y(n21) );
  MUX2XL U36 ( .D0(esfrm_wrdata[4]), .D1(memdatao[4]), .S(n2), .Y(n22) );
  MUX2XL U37 ( .D0(esfrm_wrdata[1]), .D1(memdatao[1]), .S(n2), .Y(n23) );
  MUX2XL U38 ( .D0(esfrm_wrdata[2]), .D1(memdatao[2]), .S(n2), .Y(n24) );
  MUX2XL U39 ( .D0(esfrm_wrdata[5]), .D1(memdatao[5]), .S(n2), .Y(n25) );
  INVX1 U40 ( .A(n76), .Y(n75) );
  INVX1 U41 ( .A(reset), .Y(n76) );
  BUFX3 U42 ( .A(ramdatao[0]), .Y(memdatao_comb[0]) );
  BUFX3 U43 ( .A(ramdatao[1]), .Y(memdatao_comb[1]) );
  BUFX3 U44 ( .A(ramdatao[2]), .Y(memdatao_comb[2]) );
  BUFX3 U45 ( .A(ramdatao[4]), .Y(memdatao_comb[4]) );
  BUFX3 U46 ( .A(ramdatao[5]), .Y(memdatao_comb[5]) );
  BUFX3 U47 ( .A(ramdatao[6]), .Y(memdatao_comb[6]) );
  BUFX3 U48 ( .A(ramdatao[7]), .Y(memdatao_comb[7]) );
  INVX1 U49 ( .A(n86), .Y(sfraddr[5]) );
  INVX1 U50 ( .A(n87), .Y(sfraddr[6]) );
  INVX1 U51 ( .A(sfraddr[0]), .Y(n42) );
  INVX1 U52 ( .A(n66), .Y(sfrdatao[3]) );
  INVX1 U53 ( .A(n83), .Y(ro) );
  INVX1 U54 ( .A(n60), .Y(sfrdatao[0]) );
  AO21XL U55 ( .B(sfroe_s), .C(n76), .A(esfrm_oe), .Y(sfroe) );
  INVX1 U56 ( .A(n68), .Y(sfrdatao[4]) );
  INVX1 U57 ( .A(n70), .Y(sfrdatao[5]) );
  INVX1 U58 ( .A(n72), .Y(sfrdatao[6]) );
  INVX1 U59 ( .A(n74), .Y(sfrdatao[7]) );
  INVX1 U60 ( .A(n62), .Y(sfrdatao[1]) );
  INVX1 U61 ( .A(n64), .Y(sfrdatao[2]) );
  INVX1 U62 ( .A(n87), .Y(n58) );
  NAND21XL U63 ( .B(esfrm_oe), .A(n93), .Y(sfroe_mcu51_per) );
  INVX1 U64 ( .A(n83), .Y(dbgpo[22]) );
  INVX1 U65 ( .A(n83), .Y(n81) );
  NOR21XL U66 ( .B(N19), .A(n16), .Y(N33) );
  NOR21XL U67 ( .B(N18), .A(n16), .Y(N32) );
  NOR21XL U68 ( .B(N17), .A(n16), .Y(N31) );
  NOR21XL U69 ( .B(N16), .A(n16), .Y(N30) );
  NOR21XL U70 ( .B(N15), .A(n16), .Y(N29) );
  NOR21XL U71 ( .B(N14), .A(n16), .Y(N28) );
  NOR21XL U72 ( .B(N13), .A(n6), .Y(N27) );
  NOR21XL U73 ( .B(N12), .A(n6), .Y(N26) );
  NOR21XL U74 ( .B(N11), .A(n6), .Y(N25) );
  NOR21XL U75 ( .B(N10), .A(n6), .Y(N24) );
  NOR21XL U76 ( .B(N9), .A(n6), .Y(N23) );
  NOR21XL U77 ( .B(N8), .A(n16), .Y(N22) );
  INVX1 U78 ( .A(n84), .Y(n78) );
  INVX1 U79 ( .A(n84), .Y(n77) );
  INVX1 U80 ( .A(n84), .Y(n79) );
  BUFX3 U81 ( .A(ramdatao[3]), .Y(memdatao_comb[3]) );
  BUFX3 U82 ( .A(rxd0i), .Y(dbgpo[23]) );
  MUX2IXL U83 ( .D0(esfrm_addr[4]), .D1(ramsfraddr[4]), .S(n89), .Y(n28) );
  INVX1 U84 ( .A(memdatao[3]), .Y(n88) );
  INVX1 U85 ( .A(n102), .Y(n83) );
  INVX1 U86 ( .A(n19), .Y(n60) );
  INVX1 U87 ( .A(sfroe_s), .Y(n93) );
  INVX1 U88 ( .A(n20), .Y(n72) );
  INVX1 U89 ( .A(n22), .Y(n68) );
  INVX1 U90 ( .A(n21), .Y(n74) );
  INVX1 U91 ( .A(n23), .Y(n62) );
  INVX1 U92 ( .A(n24), .Y(n64) );
  INVX1 U93 ( .A(n25), .Y(n70) );
  NOR21XL U94 ( .B(isr_irq), .A(r_hold_mcu), .Y(dbgpo[20]) );
  OR2X1 U95 ( .A(pmuintreq), .B(slp2wakeup), .Y(pmuintreq_rev) );
  OR2X1 U96 ( .A(t0_tf1), .B(t1_tf1), .Y(dbgpo[19]) );
  OR2X1 U97 ( .A(t0_tr1), .B(t1_tr1), .Y(dbgpo[18]) );
  NOR21XL U98 ( .B(N20), .A(n16), .Y(N34) );
  NOR21XL U99 ( .B(N7), .A(n6), .Y(N21) );
  NAND32X1 U100 ( .B(n11), .C(n75), .A(ien2[1]), .Y(n6) );
  INVX1 U101 ( .A(n102), .Y(n84) );
  NAND43X1 U102 ( .B(timer_1ms[8]), .C(timer_1ms[5]), .D(timer_1ms[12]), .A(
        timer_1ms[0]), .Y(n9) );
  NOR4XL U103 ( .A(n7), .B(n8), .C(n9), .D(n10), .Y(n11) );
  NAND4X1 U104 ( .A(timer_1ms[4]), .B(timer_1ms[3]), .C(timer_1ms[2]), .D(
        timer_1ms[1]), .Y(n7) );
  NAND3X1 U105 ( .A(timer_1ms[7]), .B(timer_1ms[6]), .C(timer_1ms[9]), .Y(n8)
         );
  NAND3X1 U106 ( .A(timer_1ms[11]), .B(timer_1ms[10]), .C(timer_1ms[13]), .Y(
        n10) );
  AND2X1 U107 ( .A(ien0[0]), .B(dbgpo[17]), .Y(t0_intr) );
  INVX3 U108 ( .A(esfrm_we), .Y(n91) );
  MUX2IX1 U109 ( .D0(esfrm_addr[3]), .D1(ramsfraddr[3]), .S(n2), .Y(n85) );
  INVX1 U110 ( .A(n38), .Y(n48) );
  MUX2XL U111 ( .D0(esfrm_addr[2]), .D1(ramsfraddr[2]), .S(n1), .Y(n38) );
  INVXL U112 ( .A(n48), .Y(n46) );
  INVXL U113 ( .A(n26), .Y(n44) );
  INVXL U114 ( .A(n42), .Y(n41) );
  INVX1 U115 ( .A(n90), .Y(n92) );
  INVXL U116 ( .A(n86), .Y(n103) );
  INVXL U117 ( .A(n87), .Y(n56) );
  NAND21XL U118 ( .B(n92), .A(n91), .Y(sfrwe_mcu51_per) );
  INVXL U119 ( .A(n86), .Y(n55) );
  NAND21XL U120 ( .B(isfrwait), .A(sfrwe_s), .Y(n90) );
endmodule


module mcu51_a0_DW01_inc_0 ( A, SUM );
  input [13:0] A;
  output [13:0] SUM;

  wire   [13:2] carry;

  HAD1X1 U1_1_12 ( .A(A[12]), .B(carry[12]), .CO(carry[13]), .SO(SUM[12]) );
  HAD1X1 U1_1_11 ( .A(A[11]), .B(carry[11]), .CO(carry[12]), .SO(SUM[11]) );
  HAD1X1 U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .SO(SUM[10]) );
  HAD1X1 U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .SO(SUM[9]) );
  HAD1X1 U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .SO(SUM[8]) );
  HAD1X1 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .SO(SUM[7]) );
  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  XOR2X1 U1 ( .A(carry[13]), .B(A[13]), .Y(SUM[13]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module softrstctrl_a0 ( clkcpu, resetff, newinstr, srstreq, srstflag, sfrdatai, 
        sfraddr, sfrwe );
  input [7:0] sfrdatai;
  input [6:0] sfraddr;
  input clkcpu, resetff, newinstr, sfrwe;
  output srstreq, srstflag;
  wire   srst_ff0, srst_ff1, N37, N38, N39, N40, N41, net12009, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n1, n2, n3, n4, n5, n6, n7, n8, n9;
  wire   [3:0] srst_count;

  SNPS_CLOCK_GATE_HIGH_softrstctrl_a0 clk_gate_srst_count_reg ( .CLK(clkcpu), 
        .EN(N37), .ENCLK(net12009), .TE(1'b0) );
  DFFQX1 srst_ff0_reg ( .D(n26), .C(clkcpu), .Q(srst_ff0) );
  DFFQX1 srst_ff1_reg ( .D(n24), .C(clkcpu), .Q(srst_ff1) );
  DFFQX1 srst_count_reg_1_ ( .D(N39), .C(net12009), .Q(srst_count[1]) );
  DFFQX1 srst_count_reg_0_ ( .D(N38), .C(net12009), .Q(srst_count[0]) );
  DFFQX1 srst_count_reg_3_ ( .D(N41), .C(net12009), .Q(srst_count[3]) );
  DFFQX1 srst_count_reg_2_ ( .D(N40), .C(net12009), .Q(srst_count[2]) );
  DFFQX1 srst_r_reg ( .D(n27), .C(clkcpu), .Q(srstreq) );
  DFFQX1 srstflag_reg ( .D(n25), .C(clkcpu), .Q(srstflag) );
  INVX1 U3 ( .A(n14), .Y(n2) );
  NAND42X1 U4 ( .C(sfraddr[3]), .D(n17), .A(sfraddr[0]), .B(n18), .Y(n14) );
  NAND2X1 U5 ( .A(sfraddr[2]), .B(sfraddr[1]), .Y(n17) );
  AND4X1 U6 ( .A(sfrwe), .B(sfraddr[6]), .C(sfraddr[5]), .D(sfraddr[4]), .Y(
        n18) );
  NAND2X1 U7 ( .A(sfrdatai[0]), .B(n2), .Y(n15) );
  NAND42X1 U8 ( .C(newinstr), .D(n2), .A(n9), .B(n5), .Y(n11) );
  INVX1 U9 ( .A(n12), .Y(n6) );
  NAND2X1 U10 ( .A(n9), .B(n12), .Y(N37) );
  OAI32X1 U11 ( .A(n7), .B(resetff), .C(n10), .D(n11), .E(n8), .Y(n24) );
  AOI21X1 U12 ( .B(newinstr), .C(n5), .A(n2), .Y(n10) );
  OAI22X1 U13 ( .A(n7), .B(n11), .C(resetff), .D(n15), .Y(n26) );
  NAND2X1 U14 ( .A(n12), .B(n13), .Y(n25) );
  OAI211X1 U15 ( .C(sfrdatai[0]), .D(n14), .A(n9), .B(srstflag), .Y(n13) );
  OAI33XL U16 ( .A(n16), .B(resetff), .C(n1), .D(n15), .E(resetff), .F(n8), 
        .Y(n27) );
  OAI21X1 U17 ( .B(n19), .C(n4), .A(srstreq), .Y(n16) );
  INVX1 U18 ( .A(n15), .Y(n1) );
  AOI21BBXL U19 ( .B(srst_count[1]), .C(n12), .A(N38), .Y(n21) );
  NAND2X1 U20 ( .A(srstreq), .B(n9), .Y(n12) );
  INVX1 U21 ( .A(resetff), .Y(n9) );
  OAI32X1 U22 ( .A(n19), .B(srst_count[3]), .C(n12), .D(n20), .E(n4), .Y(N41)
         );
  AOI21AX1 U23 ( .B(n6), .C(n3), .A(n21), .Y(n20) );
  NOR2X1 U24 ( .A(n12), .B(srst_count[0]), .Y(N38) );
  OAI21X1 U25 ( .B(n21), .C(n3), .A(n22), .Y(N40) );
  NAND4X1 U26 ( .A(srst_count[1]), .B(srst_count[0]), .C(n6), .D(n3), .Y(n22)
         );
  NAND3X1 U27 ( .A(srst_count[1]), .B(srst_count[0]), .C(srst_count[2]), .Y(
        n19) );
  INVX1 U28 ( .A(srst_count[3]), .Y(n4) );
  INVX1 U29 ( .A(srstreq), .Y(n5) );
  INVX1 U30 ( .A(srst_count[2]), .Y(n3) );
  NOR2X1 U31 ( .A(n23), .B(n12), .Y(N39) );
  XNOR2XL U32 ( .A(srst_count[1]), .B(srst_count[0]), .Y(n23) );
  INVX1 U33 ( .A(srst_ff0), .Y(n7) );
  INVX1 U34 ( .A(srst_ff1), .Y(n8) );
endmodule


module SNPS_CLOCK_GATE_HIGH_softrstctrl_a0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module i2c_a0 ( clk, rst, bclksel, scli, sdai, sclo, sdao, intack, si, sfrwe, 
        sfraddr, sfrdatai, i2cdat_o, i2cadr_o, i2ccon_o, i2csta_o );
  input [6:0] sfraddr;
  input [7:0] sfrdatai;
  output [7:0] i2cdat_o;
  output [7:0] i2cadr_o;
  output [7:0] i2ccon_o;
  output [7:0] i2csta_o;
  input clk, rst, bclksel, scli, sdai, intack, sfrwe;
  output sclo, sdao, si;
  wire   scli_ff, N180, sdai_ff, N181, sclo_int, wait_for_setup_r, adrcomp,
         adrcompen, nedetect, ack_bit, bsd7, pedetect, N224, N225, N226, N227,
         N232, N233, N234, sclint, ack, sdaint, bsd7_tmp, write_data_r, N296,
         N297, N298, N299, N300, N301, N302, N303, N304, N332, N333, N334,
         N335, N336, N342, N343, N344, N345, N346, N347, N348, N349, N350,
         N406, N407, N408, N409, N410, N412, N413, N414, N431, N432, N433,
         N468, N469, N470, N471, N491, N492, N493, N494, N495, busfree, N510,
         N511, rst_delay, clk_count1_ov, N653, N654, N655, N656, N657,
         clk_count2_ov, N685, N686, N687, N688, N689, N690, clkint, clkint_ff,
         N700, N746, N747, N748, N749, N1022, N1023, N1024, N1025, N1026,
         N1027, N1063, N1064, N1065, sclscl, starto_en, N1124, N1125, N1126,
         net12048, net12054, net12059, net12064, net12069, net12074, net12079,
         net12084, net12089, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
         n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n7, n8, n9, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125;
  wire   [2:0] fsmmod;
  wire   [4:0] fsmsta;
  wire   [3:0] framesync;
  wire   [2:0] fsmdet;
  wire   [2:0] setup_counter_r;
  wire   [2:0] scli_ff_reg0;
  wire   [2:0] sdai_ff_reg0;
  wire   [2:0] indelay;
  wire   [2:0] fsmsync;
  wire   [1:0] bclkcnt;
  wire   [3:0] clk_count1;
  wire   [3:0] clk_count2;

  SNPS_CLOCK_GATE_HIGH_i2c_a0_0 clk_gate_i2ccon_reg ( .CLK(clk), .EN(N224), 
        .ENCLK(net12048), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_i2c_a0_8 clk_gate_i2cdat_reg ( .CLK(clk), .EN(N296), 
        .ENCLK(net12054), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_i2c_a0_7 clk_gate_setup_counter_r_reg ( .CLK(clk), .EN(
        N332), .ENCLK(net12059), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_i2c_a0_6 clk_gate_i2cadr_reg ( .CLK(clk), .EN(N342), 
        .ENCLK(net12064), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_i2c_a0_5 clk_gate_indelay_reg ( .CLK(clk), .EN(N468), 
        .ENCLK(net12069), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_i2c_a0_4 clk_gate_framesync_reg ( .CLK(clk), .EN(N491), 
        .ENCLK(net12074), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_i2c_a0_3 clk_gate_clk_count1_reg ( .CLK(clk), .EN(N653), 
        .ENCLK(net12079), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_i2c_a0_2 clk_gate_clk_count2_reg ( .CLK(clk), .EN(N689), 
        .ENCLK(net12084), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_i2c_a0_1 clk_gate_fsmsta_reg ( .CLK(clk), .EN(N1022), 
        .ENCLK(net12089), .TE(1'b0) );
  DFFQX1 i2ccon_reg_3_ ( .D(n495), .C(clk), .Q(i2ccon_o[3]) );
  DFFQX1 scli_ff_reg ( .D(N180), .C(clk), .Q(scli_ff) );
  DFFQX1 sdai_ff_reg ( .D(N181), .C(clk), .Q(sdai_ff) );
  DFFQX1 clk_count2_ov_reg ( .D(N690), .C(clk), .Q(clk_count2_ov) );
  DFFQX1 sdai_ff_reg_reg_2_ ( .D(N433), .C(clk), .Q(sdai_ff_reg0[2]) );
  DFFQX1 clk_count2_reg_3_ ( .D(N688), .C(net12084), .Q(clk_count2[3]) );
  DFFQX1 sdai_ff_reg_reg_0_ ( .D(N431), .C(clk), .Q(sdai_ff_reg0[0]) );
  DFFQX1 sdai_ff_reg_reg_1_ ( .D(N432), .C(clk), .Q(sdai_ff_reg0[1]) );
  DFFQX1 setup_counter_r_reg_2_ ( .D(N335), .C(net12059), .Q(
        setup_counter_r[2]) );
  DFFQX1 rst_delay_reg ( .D(n24), .C(clk), .Q(rst_delay) );
  DFFQX1 clk_count1_ov_reg ( .D(n505), .C(clk), .Q(clk_count1_ov) );
  DFFQX1 bsd7_reg ( .D(n491), .C(clk), .Q(bsd7) );
  DFFQX1 ack_bit_reg ( .D(n494), .C(net12048), .Q(ack_bit) );
  DFFQX1 setup_counter_r_reg_1_ ( .D(N334), .C(net12059), .Q(
        setup_counter_r[1]) );
  DFFQX1 scli_ff_reg_reg_2_ ( .D(N414), .C(clk), .Q(scli_ff_reg0[2]) );
  DFFQX1 starto_en_reg ( .D(n490), .C(clk), .Q(starto_en) );
  DFFQX1 sclscl_reg ( .D(n59), .C(clk), .Q(sclscl) );
  DFFQX1 indelay_reg_2_ ( .D(N471), .C(net12069), .Q(indelay[2]) );
  DFFQX1 clk_count2_reg_1_ ( .D(N686), .C(net12084), .Q(clk_count2[1]) );
  DFFQX1 scli_ff_reg_reg_1_ ( .D(N413), .C(clk), .Q(scli_ff_reg0[1]) );
  DFFQX1 scli_ff_reg_reg_0_ ( .D(N412), .C(clk), .Q(scli_ff_reg0[0]) );
  DFFQX1 setup_counter_r_reg_0_ ( .D(N333), .C(net12059), .Q(
        setup_counter_r[0]) );
  DFFQX1 clk_count2_reg_0_ ( .D(N685), .C(net12084), .Q(clk_count2[0]) );
  DFFQX1 write_data_r_reg ( .D(n500), .C(clk), .Q(write_data_r) );
  DFFQX1 clk_count2_reg_2_ ( .D(N687), .C(net12084), .Q(clk_count2[2]) );
  DFFQX1 indelay_reg_1_ ( .D(N470), .C(net12069), .Q(indelay[1]) );
  DFFQX1 indelay_reg_0_ ( .D(N469), .C(net12069), .Q(indelay[0]) );
  DFFQX1 nedetect_reg ( .D(n498), .C(clk), .Q(nedetect) );
  DFFQX1 clkint_ff_reg ( .D(N700), .C(clk), .Q(clkint_ff) );
  DFFQX1 bclkcnt_reg_1_ ( .D(N511), .C(clk), .Q(bclkcnt[1]) );
  DFFQX1 bclkcnt_reg_0_ ( .D(N510), .C(clk), .Q(bclkcnt[0]) );
  DFFQX1 clk_count1_reg_2_ ( .D(N656), .C(net12079), .Q(clk_count1[2]) );
  DFFQX1 bsd7_tmp_reg ( .D(n492), .C(clk), .Q(bsd7_tmp) );
  DFFQX1 busfree_reg ( .D(n506), .C(clk), .Q(busfree) );
  DFFQX1 clk_count1_reg_3_ ( .D(N657), .C(net12079), .Q(clk_count1[3]) );
  DFFQX1 clk_count1_reg_1_ ( .D(N655), .C(net12079), .Q(clk_count1[1]) );
  DFFQX1 fsmsync_reg_1_ ( .D(N747), .C(clk), .Q(fsmsync[1]) );
  DFFQX1 clk_count1_reg_0_ ( .D(N654), .C(net12079), .Q(clk_count1[0]) );
  DFFQX1 clkint_reg ( .D(n504), .C(clk), .Q(clkint) );
  DFFQX1 adrcompen_reg ( .D(n496), .C(clk), .Q(adrcompen) );
  DFFQX1 pedetect_reg ( .D(n497), .C(clk), .Q(pedetect) );
  DFFQX1 adrcomp_reg ( .D(n501), .C(clk), .Q(adrcomp) );
  DFFQX1 fsmsync_reg_2_ ( .D(N748), .C(clk), .Q(fsmsync[2]) );
  DFFQX1 fsmsync_reg_0_ ( .D(N746), .C(clk), .Q(fsmsync[0]) );
  DFFQX1 sclint_reg ( .D(n499), .C(clk), .Q(sclint) );
  DFFQX1 fsmdet_reg_0_ ( .D(N1063), .C(clk), .Q(fsmdet[0]) );
  DFFQX1 fsmdet_reg_1_ ( .D(N1064), .C(clk), .Q(fsmdet[1]) );
  DFFQX1 fsmdet_reg_2_ ( .D(N1065), .C(clk), .Q(fsmdet[2]) );
  DFFQX1 sdaint_reg ( .D(n507), .C(clk), .Q(sdaint) );
  DFFQX1 ack_reg ( .D(n493), .C(clk), .Q(ack) );
  DFFQX1 framesync_reg_0_ ( .D(N492), .C(net12074), .Q(framesync[0]) );
  DFFQX1 framesync_reg_3_ ( .D(N495), .C(net12074), .Q(framesync[3]) );
  DFFQX1 fsmmod_reg_1_ ( .D(N1125), .C(clk), .Q(fsmmod[1]) );
  DFFQX1 fsmmod_reg_0_ ( .D(N1124), .C(clk), .Q(fsmmod[0]) );
  DFFQX1 fsmmod_reg_2_ ( .D(N1126), .C(clk), .Q(fsmmod[2]) );
  DFFQX1 fsmsta_reg_2_ ( .D(N1025), .C(net12089), .Q(fsmsta[2]) );
  DFFQX1 fsmsta_reg_3_ ( .D(N1026), .C(net12089), .Q(fsmsta[3]) );
  DFFQX1 fsmsta_reg_0_ ( .D(N1023), .C(net12089), .Q(fsmsta[0]) );
  DFFQX1 fsmsta_reg_1_ ( .D(N1024), .C(net12089), .Q(fsmsta[1]) );
  DFFQX1 framesync_reg_1_ ( .D(N493), .C(net12074), .Q(framesync[1]) );
  DFFQX1 framesync_reg_2_ ( .D(N494), .C(net12074), .Q(framesync[2]) );
  DFFQX1 fsmsta_reg_4_ ( .D(N1027), .C(net12089), .Q(fsmsta[4]) );
  DFFQX1 sclo_int_reg ( .D(N749), .C(clk), .Q(sclo_int) );
  DFFQX1 wait_for_setup_r_reg ( .D(N336), .C(clk), .Q(wait_for_setup_r) );
  DFFQX1 sdao_int_reg ( .D(n502), .C(clk), .Q(sdao) );
  DFFQX1 i2csta_reg_4_ ( .D(N410), .C(clk), .Q(i2csta_o[7]) );
  DFFQX1 i2csta_reg_3_ ( .D(N409), .C(clk), .Q(i2csta_o[6]) );
  DFFQX1 i2cdat_reg_7_ ( .D(N304), .C(net12054), .Q(i2cdat_o[7]) );
  DFFQX1 i2cadr_reg_6_ ( .D(N349), .C(net12064), .Q(i2cadr_o[6]) );
  DFFQX1 i2cadr_reg_7_ ( .D(N350), .C(net12064), .Q(i2cadr_o[7]) );
  DFFQX1 i2ccon_reg_5_ ( .D(N232), .C(net12048), .Q(i2ccon_o[5]) );
  DFFQX1 i2cadr_reg_2_ ( .D(N345), .C(net12064), .Q(i2cadr_o[2]) );
  DFFQX1 i2cdat_reg_6_ ( .D(N303), .C(net12054), .Q(i2cdat_o[6]) );
  DFFQX1 i2cdat_reg_2_ ( .D(N299), .C(net12054), .Q(i2cdat_o[2]) );
  DFFQX1 i2ccon_reg_7_ ( .D(N234), .C(net12048), .Q(i2ccon_o[7]) );
  DFFQX1 i2ccon_reg_1_ ( .D(N226), .C(net12048), .Q(i2ccon_o[1]) );
  DFFQX1 i2ccon_reg_0_ ( .D(N225), .C(net12048), .Q(i2ccon_o[0]) );
  DFFQX1 i2csta_reg_2_ ( .D(N408), .C(clk), .Q(i2csta_o[5]) );
  DFFQX1 i2csta_reg_0_ ( .D(N406), .C(clk), .Q(i2csta_o[3]) );
  DFFQX1 i2csta_reg_1_ ( .D(N407), .C(clk), .Q(i2csta_o[4]) );
  DFFQX1 i2cadr_reg_5_ ( .D(N348), .C(net12064), .Q(i2cadr_o[5]) );
  DFFQX1 i2cadr_reg_4_ ( .D(N347), .C(net12064), .Q(i2cadr_o[4]) );
  DFFQX1 i2cadr_reg_3_ ( .D(N346), .C(net12064), .Q(i2cadr_o[3]) );
  DFFQX1 i2cadr_reg_1_ ( .D(N344), .C(net12064), .Q(i2cadr_o[1]) );
  DFFQX1 i2cadr_reg_0_ ( .D(N343), .C(net12064), .Q(i2cadr_o[0]) );
  DFFQX1 i2ccon_reg_2_ ( .D(N227), .C(net12048), .Q(i2ccon_o[2]) );
  DFFQX1 i2cdat_reg_5_ ( .D(N302), .C(net12054), .Q(i2cdat_o[5]) );
  DFFQX1 i2cdat_reg_4_ ( .D(N301), .C(net12054), .Q(i2cdat_o[4]) );
  DFFQX1 i2cdat_reg_0_ ( .D(N297), .C(net12054), .Q(i2cdat_o[0]) );
  DFFQX1 i2ccon_reg_6_ ( .D(N233), .C(net12048), .Q(i2ccon_o[6]) );
  DFFQX1 i2ccon_reg_4_ ( .D(n503), .C(clk), .Q(i2ccon_o[4]) );
  DFFQX1 i2cdat_reg_3_ ( .D(N300), .C(net12054), .Q(i2cdat_o[3]) );
  DFFQX1 i2cdat_reg_1_ ( .D(N298), .C(net12054), .Q(i2cdat_o[1]) );
  INVX1 U3 ( .A(1'b1), .Y(i2csta_o[0]) );
  INVX1 U5 ( .A(1'b1), .Y(i2csta_o[1]) );
  INVX1 U7 ( .A(1'b1), .Y(i2csta_o[2]) );
  INVX1 U9 ( .A(n184), .Y(n7) );
  INVX1 U10 ( .A(si), .Y(n8) );
  NAND2X1 U11 ( .A(framesync[3]), .B(n177), .Y(n9) );
  NAND2XL U12 ( .A(sfrwe), .B(sfraddr[6]), .Y(n369) );
  AOI221XL U13 ( .A(n365), .B(n345), .C(n366), .D(n73), .E(n69), .Y(n364) );
  INVX1 U14 ( .A(N224), .Y(n32) );
  NAND2X1 U15 ( .A(n19), .B(n33), .Y(N224) );
  INVX1 U16 ( .A(n25), .Y(n19) );
  INVX1 U17 ( .A(n25), .Y(n20) );
  INVX1 U18 ( .A(n26), .Y(n21) );
  INVX1 U19 ( .A(n28), .Y(n22) );
  AOI22X1 U20 ( .A(n36), .B(n43), .C(n359), .D(n35), .Y(n163) );
  INVX1 U21 ( .A(n168), .Y(n33) );
  INVX1 U22 ( .A(n157), .Y(n36) );
  OAI21X1 U23 ( .B(n350), .C(n11), .A(n21), .Y(N343) );
  OAI21X1 U24 ( .B(n14), .C(n350), .A(n21), .Y(N346) );
  OAI21X1 U25 ( .B(n18), .C(n350), .A(n21), .Y(N350) );
  NOR2X1 U26 ( .A(n350), .B(n12), .Y(N344) );
  NOR2X1 U27 ( .A(n350), .B(n16), .Y(N348) );
  NOR2X1 U28 ( .A(n350), .B(n17), .Y(N349) );
  NOR2X1 U29 ( .A(n13), .B(n350), .Y(N345) );
  NOR2X1 U30 ( .A(n15), .B(n350), .Y(N347) );
  NAND2X1 U31 ( .A(n20), .B(n350), .Y(N342) );
  NOR2X1 U32 ( .A(n25), .B(n11), .Y(N225) );
  NOR2X1 U33 ( .A(n28), .B(n12), .Y(N226) );
  NOR2X1 U34 ( .A(n28), .B(n13), .Y(N227) );
  NOR2X1 U35 ( .A(n28), .B(n16), .Y(N232) );
  NOR2X1 U36 ( .A(n23), .B(n17), .Y(N233) );
  NOR2X1 U37 ( .A(n24), .B(n18), .Y(N234) );
  INVX1 U38 ( .A(n30), .Y(n25) );
  NAND2X1 U39 ( .A(n44), .B(n152), .Y(n359) );
  NOR2X1 U40 ( .A(n486), .B(n488), .Y(n398) );
  INVX1 U41 ( .A(n30), .Y(n26) );
  INVX1 U42 ( .A(n195), .Y(n43) );
  NOR21XL U43 ( .B(n431), .A(n69), .Y(n458) );
  INVX1 U44 ( .A(n488), .Y(n89) );
  OR2X1 U45 ( .A(n407), .B(n412), .Y(n411) );
  INVX1 U46 ( .A(n29), .Y(n24) );
  INVX1 U47 ( .A(n29), .Y(n23) );
  INVX1 U48 ( .A(n29), .Y(n27) );
  INVX1 U49 ( .A(n29), .Y(n28) );
  NOR42XL U50 ( .C(sfraddr[2]), .D(n352), .A(sfraddr[0]), .B(sfraddr[1]), .Y(
        n168) );
  NOR42XL U51 ( .C(sfraddr[1]), .D(n352), .A(sfraddr[0]), .B(sfraddr[2]), .Y(
        n157) );
  NOR42XL U52 ( .C(sfraddr[4]), .D(sfraddr[3]), .A(sfraddr[5]), .B(n369), .Y(
        n352) );
  NOR2X1 U53 ( .A(n360), .B(n361), .Y(n358) );
  AOI21X1 U54 ( .B(n360), .C(n157), .A(n361), .Y(n194) );
  INVX1 U55 ( .A(n156), .Y(n35) );
  NAND4X1 U56 ( .A(sfraddr[0]), .B(sfraddr[1]), .C(n351), .D(n352), .Y(n350)
         );
  NOR2XL U57 ( .A(sfraddr[2]), .B(n24), .Y(n351) );
  INVX1 U58 ( .A(sfrdatai[7]), .Y(n18) );
  INVX1 U59 ( .A(sfrdatai[4]), .Y(n15) );
  INVX1 U60 ( .A(sfrdatai[3]), .Y(n14) );
  INVX1 U61 ( .A(sfrdatai[5]), .Y(n16) );
  INVX1 U62 ( .A(sfrdatai[6]), .Y(n17) );
  INVX1 U63 ( .A(sfrdatai[1]), .Y(n12) );
  INVX1 U64 ( .A(sfrdatai[2]), .Y(n13) );
  INVX1 U65 ( .A(sfrdatai[0]), .Y(n11) );
  OR2X1 U66 ( .A(sdai), .B(n27), .Y(N181) );
  INVX1 U67 ( .A(n150), .Y(n44) );
  INVX1 U68 ( .A(rst), .Y(n30) );
  NAND2X1 U69 ( .A(n363), .B(n65), .Y(n152) );
  INVX1 U70 ( .A(n181), .Y(n91) );
  NOR32XL U71 ( .B(n489), .C(n488), .A(n486), .Y(n402) );
  NAND2X1 U72 ( .A(n363), .B(n364), .Y(n195) );
  NAND4X1 U73 ( .A(n442), .B(n434), .C(n438), .D(n444), .Y(n465) );
  NAND3X1 U74 ( .A(n172), .B(n20), .C(n173), .Y(n486) );
  NAND2X1 U75 ( .A(n475), .B(n73), .Y(n457) );
  NOR2X1 U76 ( .A(n468), .B(n478), .Y(n442) );
  AOI21X1 U77 ( .B(n423), .C(n432), .A(n112), .Y(n456) );
  INVX1 U78 ( .A(n364), .Y(n65) );
  INVX1 U79 ( .A(n203), .Y(n67) );
  INVX1 U80 ( .A(n404), .Y(n69) );
  INVX1 U81 ( .A(n183), .Y(n56) );
  NOR2X1 U82 ( .A(n90), .B(n334), .Y(n488) );
  NAND2X1 U83 ( .A(n78), .B(n365), .Y(n263) );
  NAND2X1 U84 ( .A(n482), .B(n73), .Y(n340) );
  NAND2X1 U85 ( .A(n482), .B(n70), .Y(n431) );
  INVX1 U86 ( .A(n365), .Y(n63) );
  INVX1 U87 ( .A(n236), .Y(n55) );
  NAND2X1 U88 ( .A(n434), .B(n435), .Y(n407) );
  NAND3X1 U89 ( .A(n428), .B(n340), .C(n429), .Y(n409) );
  NAND3X1 U90 ( .A(n203), .B(n443), .C(n444), .Y(n440) );
  NAND2X1 U91 ( .A(n431), .B(n432), .Y(n412) );
  INVX1 U92 ( .A(n336), .Y(n116) );
  INVX1 U93 ( .A(rst), .Y(n29) );
  OR2X1 U94 ( .A(n268), .B(n119), .Y(n273) );
  INVX1 U95 ( .A(n334), .Y(n92) );
  INVX1 U96 ( .A(n249), .Y(n103) );
  INVX1 U97 ( .A(n320), .Y(n84) );
  INVX1 U98 ( .A(n246), .Y(n40) );
  INVX1 U99 ( .A(n281), .Y(n118) );
  OAI32X1 U100 ( .A(n33), .B(n26), .C(n31), .D(n109), .E(n230), .Y(n503) );
  INVX1 U101 ( .A(n230), .Y(n31) );
  OAI221X1 U102 ( .A(n168), .B(n231), .C(n33), .D(n15), .E(n22), .Y(n230) );
  AOI21X1 U103 ( .B(n107), .C(n232), .A(n233), .Y(n231) );
  OAI21X1 U104 ( .B(n154), .C(n98), .A(n155), .Y(n492) );
  GEN2XL U105 ( .D(n156), .E(n18), .C(n44), .B(n22), .A(n34), .Y(n155) );
  INVX1 U106 ( .A(n154), .Y(n34) );
  OAI21BBX1 U107 ( .A(n148), .B(n157), .C(n145), .Y(n154) );
  NAND2X1 U108 ( .A(n36), .B(n8), .Y(n156) );
  ENOX1 U109 ( .A(n36), .B(n195), .C(n359), .D(n149), .Y(n361) );
  OAI22X1 U110 ( .A(n358), .B(n14), .C(n163), .D(n97), .Y(N300) );
  OAI22X1 U111 ( .A(n358), .B(n13), .C(n163), .D(n96), .Y(N299) );
  OAI22X1 U112 ( .A(n358), .B(n12), .C(n163), .D(n81), .Y(N298) );
  OAI22X1 U113 ( .A(n358), .B(n11), .C(n163), .D(n95), .Y(N297) );
  AOI22X1 U114 ( .A(n148), .B(n36), .C(n149), .D(n150), .Y(n147) );
  OAI211X1 U115 ( .C(n362), .D(n87), .A(n194), .B(n21), .Y(N296) );
  AOI21X1 U116 ( .B(n35), .C(n359), .A(n43), .Y(n362) );
  OAI21X1 U117 ( .B(n160), .C(n95), .A(n161), .Y(n493) );
  OAI21BBX1 U118 ( .A(n52), .B(n162), .C(n160), .Y(n161) );
  OAI21X1 U119 ( .B(n163), .C(n87), .A(n162), .Y(n160) );
  NOR2X1 U120 ( .A(n24), .B(n148), .Y(n162) );
  OR2X1 U121 ( .A(scli), .B(n27), .Y(N180) );
  NOR32XL U122 ( .B(n91), .C(n225), .A(n45), .Y(n363) );
  INVX1 U123 ( .A(n453), .Y(n46) );
  OAI221X1 U124 ( .A(n433), .B(n435), .C(n111), .D(n340), .E(n454), .Y(n453)
         );
  AOI211X1 U125 ( .C(n51), .D(n455), .A(n71), .B(n456), .Y(n454) );
  INVX1 U126 ( .A(n457), .Y(n71) );
  NOR3XL U127 ( .A(n45), .B(n225), .C(n181), .Y(n150) );
  NAND2X1 U128 ( .A(n483), .B(n73), .Y(n423) );
  INVX1 U129 ( .A(n184), .Y(n112) );
  NAND2X1 U130 ( .A(n19), .B(n182), .Y(n181) );
  OAI2B11X1 U131 ( .D(n359), .C(n83), .A(n158), .B(n196), .Y(n360) );
  NAND2X1 U132 ( .A(n480), .B(n70), .Y(n427) );
  OAI221X1 U133 ( .A(n112), .B(n390), .C(n9), .D(n427), .E(n423), .Y(n455) );
  OAI211X1 U134 ( .C(n82), .D(n413), .A(n447), .B(n448), .Y(N1024) );
  AOI31X1 U135 ( .A(n205), .B(n95), .C(n402), .D(n54), .Y(n448) );
  OAI31XL U136 ( .A(n449), .B(n450), .C(n451), .D(n400), .Y(n447) );
  INVX1 U137 ( .A(n414), .Y(n54) );
  NOR2X1 U138 ( .A(n83), .B(n44), .Y(n148) );
  OAI211X1 U139 ( .C(n125), .D(n432), .A(n46), .B(n50), .Y(n451) );
  INVX1 U140 ( .A(n452), .Y(n50) );
  NAND31X1 U141 ( .C(n174), .A(n398), .B(n179), .Y(n414) );
  NOR21XL U142 ( .B(n366), .A(n77), .Y(n482) );
  NAND31X1 U143 ( .C(n330), .A(n66), .B(n366), .Y(n432) );
  AOI22X1 U144 ( .A(n70), .B(n475), .C(n475), .D(n481), .Y(n434) );
  AND2X1 U145 ( .A(n368), .B(n73), .Y(n478) );
  AND2X1 U146 ( .A(n368), .B(n348), .Y(n468) );
  INVX1 U147 ( .A(n264), .Y(n73) );
  OAI21X1 U148 ( .B(n200), .C(n112), .A(n65), .Y(n224) );
  NAND2X1 U149 ( .A(n348), .B(n483), .Y(n203) );
  NOR2X1 U150 ( .A(n109), .B(n202), .Y(n183) );
  NAND2X1 U151 ( .A(n70), .B(n479), .Y(n404) );
  AND2X1 U152 ( .A(n224), .B(n218), .Y(n223) );
  AOI21X1 U153 ( .B(n95), .C(n402), .A(n28), .Y(n417) );
  INVX1 U154 ( .A(n331), .Y(n70) );
  NOR2X1 U155 ( .A(n341), .B(n75), .Y(n475) );
  NAND41X1 U156 ( .D(n476), .A(n403), .B(n443), .C(n477), .Y(n452) );
  NAND3X1 U157 ( .A(n184), .B(n408), .C(n478), .Y(n477) );
  OAI22X1 U158 ( .A(n429), .B(n446), .C(n428), .D(n111), .Y(n476) );
  OAI211X1 U159 ( .C(n111), .D(n429), .A(n46), .B(n445), .Y(n439) );
  OA222X1 U160 ( .A(n431), .B(n112), .C(n446), .D(n428), .E(n433), .F(n434), 
        .Y(n445) );
  OAI22AX1 U161 ( .D(n216), .C(n217), .A(n216), .B(n125), .Y(n502) );
  AOI211X1 U162 ( .C(n218), .D(n219), .A(n220), .B(n42), .Y(n217) );
  NAND3X1 U163 ( .A(n221), .B(n218), .C(n226), .Y(n216) );
  INVX1 U164 ( .A(n221), .Y(n42) );
  AOI211X1 U165 ( .C(n473), .D(n425), .A(n452), .B(n410), .Y(n472) );
  NAND4X1 U166 ( .A(n458), .B(n427), .C(n423), .D(n340), .Y(n473) );
  NAND2X1 U167 ( .A(n368), .B(n74), .Y(n390) );
  NAND3X1 U168 ( .A(n381), .B(n382), .C(n227), .Y(n202) );
  NOR2X1 U169 ( .A(n229), .B(n282), .Y(n381) );
  NAND2X1 U170 ( .A(n481), .B(n483), .Y(n444) );
  NAND2X1 U171 ( .A(n483), .B(n70), .Y(n438) );
  NAND2X1 U172 ( .A(n45), .B(n19), .Y(n196) );
  NAND2X1 U173 ( .A(n480), .B(n73), .Y(n428) );
  NAND2X1 U174 ( .A(n481), .B(n482), .Y(n429) );
  NAND2X1 U175 ( .A(n112), .B(n125), .Y(n446) );
  INVX1 U176 ( .A(n425), .Y(n111) );
  NAND42X1 U177 ( .C(n402), .D(n400), .A(n414), .B(n485), .Y(N1022) );
  NOR21XL U178 ( .B(n413), .A(n486), .Y(n485) );
  NOR2X1 U179 ( .A(n310), .B(n23), .Y(n236) );
  NOR4XL U180 ( .A(n486), .B(n89), .C(n87), .D(n489), .Y(n400) );
  NOR2X1 U181 ( .A(n93), .B(n395), .Y(n334) );
  NAND3X1 U182 ( .A(n121), .B(n20), .C(n260), .Y(n336) );
  NAND2X1 U183 ( .A(n75), .B(n66), .Y(n365) );
  AOI221XL U184 ( .A(n407), .B(n408), .C(n111), .D(n409), .E(n410), .Y(n406)
         );
  AOI22AXL U185 ( .A(n433), .B(n407), .D(n427), .C(n408), .Y(n418) );
  NOR3XL U186 ( .A(n390), .B(n95), .C(n9), .Y(n430) );
  NOR3XL U187 ( .A(n87), .B(n67), .C(n426), .Y(n489) );
  NOR2X1 U188 ( .A(n100), .B(n62), .Y(n282) );
  OAI221X1 U189 ( .A(n252), .B(n181), .C(n115), .D(n181), .E(n22), .Y(n506) );
  AOI21BX1 U190 ( .C(n253), .B(n232), .A(n233), .Y(n252) );
  OAI31XL U191 ( .A(n353), .B(n355), .C(n99), .D(n354), .Y(N335) );
  NAND3X1 U192 ( .A(n90), .B(n58), .C(n282), .Y(n173) );
  INVX1 U193 ( .A(n182), .Y(n90) );
  NAND2X1 U194 ( .A(n475), .B(n348), .Y(n435) );
  NAND2X1 U195 ( .A(n73), .B(n479), .Y(n403) );
  NOR2X1 U196 ( .A(n297), .B(n291), .Y(N687) );
  XNOR2XL U197 ( .A(n293), .B(n106), .Y(n297) );
  NAND2X1 U198 ( .A(n383), .B(n90), .Y(n172) );
  NAND2X1 U199 ( .A(n430), .B(n52), .Y(n443) );
  INVX1 U200 ( .A(n349), .Y(n78) );
  INVX1 U201 ( .A(n142), .Y(n61) );
  NAND2X1 U202 ( .A(n353), .B(n354), .Y(N336) );
  NAND2X1 U203 ( .A(n236), .B(n108), .Y(N700) );
  NAND2X1 U204 ( .A(n236), .B(n105), .Y(N689) );
  INVX1 U205 ( .A(n408), .Y(n51) );
  INVX1 U206 ( .A(n205), .Y(n80) );
  INVX1 U207 ( .A(n341), .Y(n76) );
  OAI21X1 U208 ( .B(n309), .C(n102), .A(n103), .Y(n245) );
  AOI211X1 U209 ( .C(n82), .D(n228), .A(n229), .B(n45), .Y(n221) );
  AND4X1 U210 ( .A(n107), .B(n228), .C(n83), .D(n109), .Y(n378) );
  INVX1 U211 ( .A(n178), .Y(n113) );
  NOR2X1 U212 ( .A(n104), .B(n309), .Y(n249) );
  NOR2X1 U213 ( .A(n328), .B(n7), .Y(n320) );
  NAND2X1 U214 ( .A(n289), .B(n120), .Y(n281) );
  NOR2X1 U215 ( .A(n83), .B(n23), .Y(n338) );
  OAI222XL U216 ( .A(n240), .B(n241), .C(n242), .D(n243), .E(n101), .F(n244), 
        .Y(n239) );
  INVX1 U217 ( .A(n245), .Y(n101) );
  NAND3X1 U218 ( .A(n47), .B(n41), .C(n48), .Y(n246) );
  NOR2X1 U219 ( .A(n102), .B(n104), .Y(n302) );
  OAI21X1 U220 ( .B(n78), .C(n346), .A(n338), .Y(N408) );
  XNOR2XL U221 ( .A(n264), .B(n75), .Y(n346) );
  OAI21X1 U222 ( .B(n323), .C(n84), .A(n91), .Y(N494) );
  XNOR2XL U223 ( .A(n322), .B(n114), .Y(n323) );
  INVX1 U224 ( .A(n305), .Y(n38) );
  OAI211X1 U225 ( .C(n244), .D(n245), .A(n306), .B(n307), .Y(n305) );
  AOI211X1 U226 ( .C(n250), .D(n103), .A(n251), .B(n40), .Y(n307) );
  AOI22AXL U227 ( .A(n39), .B(n243), .D(n241), .C(n240), .Y(n306) );
  NOR2X1 U228 ( .A(n280), .B(n283), .Y(n268) );
  AOI21X1 U229 ( .B(n264), .C(n75), .A(n77), .Y(n262) );
  NAND2X1 U230 ( .A(n20), .B(n313), .Y(n317) );
  OAI211X1 U231 ( .C(n77), .D(n342), .A(n338), .B(n343), .Y(N409) );
  AOI22AXL U232 ( .A(n344), .B(n77), .D(n344), .C(n345), .Y(n343) );
  NOR2X1 U233 ( .A(n264), .B(n75), .Y(n344) );
  OAI21AX1 U234 ( .B(n86), .C(n190), .A(n186), .Y(n499) );
  OR2X1 U235 ( .A(n228), .B(n27), .Y(n267) );
  NAND4X1 U236 ( .A(n327), .B(n91), .C(n113), .D(n328), .Y(N491) );
  NAND2X1 U237 ( .A(n20), .B(n187), .Y(n186) );
  INVX1 U238 ( .A(n388), .Y(n107) );
  NAND2X1 U239 ( .A(n338), .B(n347), .Y(N407) );
  OAI21X1 U240 ( .B(n348), .C(n70), .A(n349), .Y(n347) );
  NAND2X1 U241 ( .A(n116), .B(n271), .Y(N468) );
  INVX1 U242 ( .A(n285), .Y(n119) );
  INVX1 U243 ( .A(n242), .Y(n39) );
  INVX1 U244 ( .A(n313), .Y(n37) );
  NOR21XL U245 ( .B(n260), .A(n271), .Y(n278) );
  NOR2X1 U246 ( .A(n93), .B(n94), .Y(n394) );
  NOR2X1 U247 ( .A(n120), .B(n117), .Y(n260) );
  NOR2X1 U248 ( .A(n121), .B(n120), .Y(n270) );
  NAND2X1 U249 ( .A(n63), .B(n74), .Y(n342) );
  INVX1 U250 ( .A(n190), .Y(n49) );
  NAND2X1 U251 ( .A(n388), .B(n280), .Y(n377) );
  NAND2X1 U252 ( .A(n283), .B(n285), .Y(n284) );
  INVX1 U253 ( .A(n382), .Y(n57) );
  ENOX1 U254 ( .A(n166), .B(n167), .C(i2ccon_o[3]), .D(n166), .Y(n495) );
  AOI32X1 U255 ( .A(n168), .B(n20), .C(sfrdatai[3]), .D(n169), .E(n32), .Y(
        n167) );
  NOR32XL U256 ( .B(n170), .C(n20), .A(n169), .Y(n166) );
  AOI31X1 U257 ( .A(n171), .B(n172), .C(n173), .D(n45), .Y(n169) );
  AO22AXL U258 ( .A(n143), .B(n144), .C(bsd7), .D(n144), .Y(n491) );
  OAI211X1 U259 ( .C(n151), .D(n44), .A(n21), .B(n146), .Y(n143) );
  NAND3X1 U260 ( .A(n145), .B(n146), .C(n147), .Y(n144) );
  NOR21XL U261 ( .B(n152), .A(n43), .Y(n146) );
  OAI22AX1 U262 ( .D(i2cdat_o[6]), .C(n163), .A(n358), .B(n18), .Y(N304) );
  OAI22AX1 U263 ( .D(i2cdat_o[5]), .C(n163), .A(n358), .B(n17), .Y(N303) );
  OAI22AX1 U264 ( .D(i2cdat_o[4]), .C(n163), .A(n358), .B(n16), .Y(N302) );
  OAI22AX1 U265 ( .D(i2cdat_o[3]), .C(n163), .A(n358), .B(n15), .Y(N301) );
  AOI221XL U266 ( .A(sfrdatai[7]), .B(n149), .C(i2cdat_o[7]), .D(n35), .E(n153), .Y(n151) );
  AOI21X1 U267 ( .B(n86), .C(n98), .A(n83), .Y(n153) );
  OAI21X1 U268 ( .B(n192), .C(n193), .A(n194), .Y(n500) );
  NAND4X1 U269 ( .A(write_data_r), .B(n168), .C(n195), .D(n44), .Y(n193) );
  NAND4X1 U270 ( .A(n158), .B(n196), .C(n156), .D(n19), .Y(n192) );
  AOI22X1 U271 ( .A(intack), .B(n33), .C(n168), .D(n14), .Y(n170) );
  NOR2X1 U272 ( .A(n36), .B(i2ccon_o[3]), .Y(n149) );
  NOR32XL U273 ( .B(n158), .C(n159), .A(n27), .Y(n145) );
  NAND4X1 U274 ( .A(nedetect), .B(n35), .C(n150), .D(n87), .Y(n159) );
  OAI21BX1 U275 ( .C(ack_bit), .B(n164), .A(n165), .Y(n494) );
  OAI21X1 U276 ( .B(sfrdatai[2]), .C(n28), .A(n164), .Y(n165) );
  OAI31XL U277 ( .A(n33), .B(n83), .C(n152), .D(n21), .Y(n164) );
  AND2X1 U278 ( .A(sclo_int), .B(n85), .Y(sclo) );
  INVX1 U279 ( .A(wait_for_setup_r), .Y(n85) );
  NOR21XL U280 ( .B(n366), .A(fsmsta[3]), .Y(n483) );
  NOR21XL U281 ( .B(n345), .A(fsmsta[2]), .Y(n480) );
  NAND2X1 U282 ( .A(framesync[3]), .B(n177), .Y(n184) );
  NOR3XL U283 ( .A(framesync[1]), .B(framesync[2]), .C(framesync[0]), .Y(n177)
         );
  NOR2X1 U284 ( .A(n75), .B(fsmsta[4]), .Y(n366) );
  NOR2X1 U285 ( .A(n77), .B(fsmsta[4]), .Y(n345) );
  GEN2XL U286 ( .D(framesync[3]), .E(n222), .C(bsd7), .B(n223), .A(n24), .Y(
        n220) );
  NAND2X1 U287 ( .A(fsmsta[4]), .B(n77), .Y(n341) );
  INVX1 U288 ( .A(fsmsta[3]), .Y(n77) );
  INVX1 U289 ( .A(fsmsta[1]), .Y(n74) );
  NAND2X1 U290 ( .A(fsmsta[0]), .B(fsmsta[1]), .Y(n264) );
  INVX1 U291 ( .A(fsmsta[2]), .Y(n75) );
  NAND2X1 U292 ( .A(sdao), .B(n112), .Y(n425) );
  NOR3XL U293 ( .A(fsmmod[1]), .B(fsmmod[2]), .C(n58), .Y(n383) );
  NOR3XL U294 ( .A(fsmsta[3]), .B(fsmsta[4]), .C(fsmsta[2]), .Y(n368) );
  NOR3XL U295 ( .A(n58), .B(fsmmod[2]), .C(n100), .Y(n229) );
  NAND2X1 U296 ( .A(fsmsta[0]), .B(n74), .Y(n331) );
  NOR2X1 U297 ( .A(n74), .B(fsmsta[0]), .Y(n348) );
  OAI222XL U298 ( .A(n458), .B(n425), .C(n459), .D(n203), .E(n460), .F(n9), 
        .Y(n450) );
  AOI31X1 U299 ( .A(n80), .B(n95), .C(i2cadr_o[0]), .D(n426), .Y(n459) );
  AOI22BXL U300 ( .B(n434), .A(n461), .D(n390), .C(n95), .Y(n460) );
  OR2X1 U301 ( .A(i2ccon_o[2]), .B(sdaint), .Y(n461) );
  AOI21X1 U302 ( .B(n58), .C(fsmmod[2]), .A(n383), .Y(n227) );
  NOR2X1 U303 ( .A(fsmsta[1]), .B(fsmsta[0]), .Y(n481) );
  NOR2X1 U304 ( .A(n341), .B(fsmsta[2]), .Y(n479) );
  NOR3XL U305 ( .A(i2ccon_o[2]), .B(sdaint), .C(n184), .Y(n433) );
  OAI211X1 U306 ( .C(n426), .D(n474), .A(n457), .B(n263), .Y(n410) );
  NAND2X1 U307 ( .A(n67), .B(ack), .Y(n474) );
  INVX1 U308 ( .A(fsmmod[0]), .Y(n58) );
  AOI211X1 U309 ( .C(n200), .D(nedetect), .A(n27), .B(n223), .Y(n226) );
  OAI21BX1 U310 ( .C(n400), .B(n436), .A(n437), .Y(N1025) );
  OAI21X1 U311 ( .B(n80), .C(ack), .A(n402), .Y(n437) );
  NOR41XL U312 ( .D(n438), .A(n439), .B(n440), .C(n441), .Y(n436) );
  AOI21X1 U313 ( .B(n408), .C(n9), .A(n442), .Y(n441) );
  INVX1 U314 ( .A(fsmmod[1]), .Y(n100) );
  NAND3X1 U315 ( .A(n90), .B(n21), .C(i2ccon_o[6]), .Y(n158) );
  ENOX1 U316 ( .A(ack_bit), .B(n224), .C(n224), .D(n225), .Y(n219) );
  OAI211X1 U317 ( .C(ack), .D(n390), .A(n435), .B(n68), .Y(n484) );
  INVX1 U318 ( .A(n465), .Y(n68) );
  OAI211X1 U319 ( .C(n425), .D(n427), .A(n463), .B(n464), .Y(n449) );
  AOI32X1 U320 ( .A(n63), .B(fsmsta[1]), .C(n78), .D(n468), .E(n184), .Y(n463)
         );
  AOI31X1 U321 ( .A(n465), .B(n184), .C(n51), .D(n466), .Y(n464) );
  OAI21X1 U322 ( .B(n125), .C(n423), .A(n467), .Y(n466) );
  OAI211X1 U323 ( .C(adrcomp), .D(n413), .A(n414), .B(n415), .Y(N1026) );
  AOI21AX1 U324 ( .B(n400), .C(n416), .A(n417), .Y(n415) );
  NAND4X1 U325 ( .A(n418), .B(n419), .C(n420), .D(n421), .Y(n416) );
  AOI22X1 U326 ( .A(n430), .B(sdaint), .C(n412), .D(n184), .Y(n419) );
  NAND3X1 U327 ( .A(n92), .B(n56), .C(i2ccon_o[6]), .Y(n233) );
  NAND2X1 U328 ( .A(fsmsta[3]), .B(fsmsta[1]), .Y(n330) );
  NAND4X1 U329 ( .A(n417), .B(n173), .C(n469), .D(n413), .Y(N1023) );
  NAND2X1 U330 ( .A(n400), .B(n470), .Y(n469) );
  OAI211X1 U331 ( .C(n446), .D(n432), .A(n471), .B(n472), .Y(n470) );
  AOI33X1 U332 ( .A(n9), .B(n408), .C(n70), .D(sdaint), .E(n484), .F(n112), 
        .Y(n471) );
  NOR21XL U333 ( .B(framesync[3]), .A(n222), .Y(n178) );
  NAND31X1 U334 ( .C(framesync[1]), .A(n114), .B(framesync[0]), .Y(n222) );
  AO22AXL U335 ( .A(n355), .B(n99), .C(n188), .D(n357), .Y(n353) );
  NOR2X1 U336 ( .A(write_data_r), .B(n23), .Y(n357) );
  GEN2XL U337 ( .D(framesync[3]), .E(n319), .C(n200), .B(n320), .A(n321), .Y(
        N495) );
  OR2X1 U338 ( .A(n322), .B(n114), .Y(n319) );
  XNOR2XL U339 ( .A(i2cdat_o[6]), .B(i2cadr_o[7]), .Y(n215) );
  OA22X1 U340 ( .A(n174), .B(n175), .C(n82), .D(n176), .Y(n171) );
  OAI21X1 U341 ( .B(n177), .C(n178), .A(n89), .Y(n176) );
  AOI22X1 U342 ( .A(n112), .B(pedetect), .C(n179), .D(n89), .Y(n175) );
  OAI21X1 U343 ( .B(n487), .C(n375), .A(n398), .Y(n413) );
  NOR32XL U344 ( .B(n177), .C(n83), .A(framesync[3]), .Y(n487) );
  XNOR2XL U345 ( .A(i2cdat_o[1]), .B(i2cadr_o[2]), .Y(n209) );
  XNOR2XL U346 ( .A(i2cdat_o[4]), .B(i2cadr_o[5]), .Y(n210) );
  XNOR2XL U347 ( .A(i2cdat_o[0]), .B(i2cadr_o[1]), .Y(n211) );
  NAND21X1 U348 ( .B(scli_ff_reg0[1]), .A(n19), .Y(N414) );
  NAND21X1 U349 ( .B(scli_ff_reg0[0]), .A(n19), .Y(N413) );
  NAND32X1 U350 ( .B(n398), .C(n26), .A(n399), .Y(N1027) );
  AOI22X1 U351 ( .A(n400), .B(n401), .C(n402), .D(ack), .Y(n399) );
  NAND4X1 U352 ( .A(n403), .B(n404), .C(n405), .D(n406), .Y(n401) );
  AOI22X1 U353 ( .A(n63), .B(fsmsta[4]), .C(n112), .D(n411), .Y(n405) );
  OAI21X1 U354 ( .B(framesync[3]), .C(n177), .A(n184), .Y(n179) );
  NAND2X1 U355 ( .A(sdao), .B(n52), .Y(n408) );
  INVX1 U356 ( .A(sdaint), .Y(n52) );
  NAND4X1 U357 ( .A(n96), .B(n97), .C(n81), .D(n462), .Y(n205) );
  NOR4XL U358 ( .A(i2cdat_o[6]), .B(i2cdat_o[5]), .C(i2cdat_o[4]), .D(
        i2cdat_o[3]), .Y(n462) );
  AND2X1 U359 ( .A(i2ccon_o[5]), .B(n390), .Y(n333) );
  AOI21AX1 U360 ( .B(adrcomp), .C(adrcompen), .A(n227), .Y(n218) );
  NAND3X1 U361 ( .A(fsmdet[0]), .B(n93), .C(fsmdet[1]), .Y(n182) );
  INVX1 U362 ( .A(fsmsta[0]), .Y(n66) );
  AOI221XL U363 ( .A(n63), .B(fsmsta[3]), .C(n422), .D(n72), .E(n64), .Y(n421)
         );
  INVX1 U364 ( .A(n263), .Y(n64) );
  NOR2X1 U365 ( .A(n51), .B(n9), .Y(n422) );
  INVX1 U366 ( .A(n423), .Y(n72) );
  NAND3X1 U367 ( .A(n58), .B(n62), .C(fsmmod[1]), .Y(n382) );
  NOR3XL U368 ( .A(n322), .B(framesync[3]), .C(n114), .Y(n200) );
  AOI211X1 U369 ( .C(n202), .D(n203), .A(n204), .B(n88), .Y(n201) );
  OAI21X1 U370 ( .B(n95), .C(n205), .A(n206), .Y(n204) );
  ENOX1 U371 ( .A(n207), .B(n208), .C(n80), .D(i2cadr_o[0]), .Y(n206) );
  NAND3X1 U372 ( .A(n209), .B(n210), .C(n211), .Y(n208) );
  NAND2X1 U373 ( .A(fsmsta[3]), .B(fsmsta[4]), .Y(n349) );
  AOI31X1 U374 ( .A(fsmsta[2]), .B(n77), .C(n367), .D(n368), .Y(n225) );
  OAI21X1 U375 ( .B(n79), .C(fsmsta[0]), .A(fsmsta[1]), .Y(n367) );
  NAND3X1 U376 ( .A(fsmmod[0]), .B(n100), .C(fsmmod[2]), .Y(n142) );
  INVX1 U377 ( .A(ack), .Y(n95) );
  NAND2X1 U378 ( .A(clk_count1_ov), .B(n236), .Y(n291) );
  INVX1 U379 ( .A(fsmsta[4]), .Y(n79) );
  OAI32X1 U380 ( .A(n87), .B(n185), .C(n186), .D(sclint), .E(n187), .Y(n497)
         );
  OAI32X1 U381 ( .A(n55), .B(n38), .C(n303), .D(n26), .E(n285), .Y(N656) );
  XNOR2XL U382 ( .A(n302), .B(clk_count1[2]), .Y(n303) );
  EORX1 U383 ( .A(n424), .B(n425), .C(n426), .D(ack), .Y(n420) );
  NAND21X1 U384 ( .B(n409), .A(n427), .Y(n424) );
  INVX1 U385 ( .A(sdao), .Y(n125) );
  NOR3XL U386 ( .A(fsmmod[0]), .B(fsmmod[1]), .C(n62), .Y(n232) );
  NAND2X1 U387 ( .A(sclint), .B(n19), .Y(n188) );
  AOI31X1 U388 ( .A(scli_ff_reg0[2]), .B(N414), .C(N413), .D(n190), .Y(n185)
         );
  OAI211X1 U389 ( .C(n325), .D(n326), .A(n91), .B(n327), .Y(n321) );
  AOI21BBXL U390 ( .B(n328), .C(n9), .A(n329), .Y(n326) );
  NOR3XL U391 ( .A(n333), .B(i2ccon_o[4]), .C(i2ccon_o[3]), .Y(n325) );
  AOI31X1 U392 ( .A(n330), .B(n331), .C(n332), .D(n113), .Y(n329) );
  INVX1 U393 ( .A(fsmmod[2]), .Y(n62) );
  OAI21X1 U394 ( .B(clk_count2[0]), .C(n55), .A(n299), .Y(N685) );
  NAND4X1 U395 ( .A(fsmsync[2]), .B(n117), .C(n120), .D(n19), .Y(n299) );
  OAI21X1 U396 ( .B(n49), .C(n188), .A(n189), .Y(n498) );
  NAND42X1 U397 ( .C(n185), .D(n190), .A(nedetect), .B(n19), .Y(n189) );
  OAI21X1 U398 ( .B(n108), .C(n234), .A(n235), .Y(n504) );
  OAI21X1 U399 ( .B(n55), .C(n108), .A(n234), .Y(n235) );
  NAND21X1 U400 ( .B(clk_count2_ov), .A(n236), .Y(n234) );
  OAI31XL U401 ( .A(n53), .B(n27), .C(n105), .D(n237), .Y(n505) );
  OAI211X1 U402 ( .C(n238), .D(n239), .A(n53), .B(n236), .Y(n237) );
  INVX1 U403 ( .A(rst_delay), .Y(n53) );
  OAI31XL U404 ( .A(n246), .B(n103), .C(n102), .D(n247), .Y(n238) );
  OAI21X1 U405 ( .B(rst_delay), .C(n311), .A(n21), .Y(N653) );
  NOR4XL U406 ( .A(n312), .B(n310), .C(n37), .D(n39), .Y(n311) );
  NAND42X1 U407 ( .C(n250), .D(n40), .A(n241), .B(n244), .Y(n312) );
  INVX1 U408 ( .A(fsmdet[2]), .Y(n93) );
  GEN2XL U409 ( .D(n116), .E(n123), .C(N469), .B(indelay[2]), .A(n335), .Y(
        N471) );
  NOR4XL U410 ( .A(indelay[2]), .B(n123), .C(n336), .D(n122), .Y(n335) );
  INVX1 U411 ( .A(indelay[1]), .Y(n123) );
  INVX1 U412 ( .A(indelay[0]), .Y(n122) );
  INVX1 U413 ( .A(fsmdet[1]), .Y(n94) );
  NAND3X1 U414 ( .A(n112), .B(adrcomp), .C(adrcompen), .Y(n426) );
  NAND3X1 U415 ( .A(n92), .B(n56), .C(n314), .Y(n310) );
  AOI22AXL U416 ( .A(n315), .B(n86), .D(n289), .C(n120), .Y(n314) );
  ENOX1 U417 ( .A(n61), .B(n115), .C(sclo_int), .D(n232), .Y(n315) );
  NAND2X1 U418 ( .A(fsmdet[0]), .B(n94), .Y(n395) );
  OAI2B11X1 U419 ( .D(write_data_r), .C(sclint), .A(n353), .B(n21), .Y(N332)
         );
  NOR3XL U420 ( .A(n55), .B(n38), .C(n300), .Y(N657) );
  XNOR2XL U421 ( .A(clk_count1[3]), .B(n301), .Y(n300) );
  AND2X1 U422 ( .A(clk_count1[2]), .B(n302), .Y(n301) );
  NOR3XL U423 ( .A(n55), .B(n38), .C(n304), .Y(N655) );
  XNOR2XL U424 ( .A(clk_count1[1]), .B(clk_count1[0]), .Y(n304) );
  NOR3XL U425 ( .A(n55), .B(clk_count1[0]), .C(n38), .Y(N654) );
  OAI211X1 U426 ( .C(n345), .D(n76), .A(fsmsta[1]), .B(n63), .Y(n467) );
  NAND2X1 U427 ( .A(framesync[1]), .B(framesync[0]), .Y(n322) );
  NOR2X1 U428 ( .A(n202), .B(adrcomp), .Y(n174) );
  NOR2X1 U429 ( .A(n336), .B(indelay[0]), .Y(N469) );
  OAI21AX1 U430 ( .B(framesync[0]), .C(n84), .A(n321), .Y(N492) );
  NOR2X1 U431 ( .A(n356), .B(n353), .Y(N334) );
  AOI21X1 U432 ( .B(setup_counter_r[1]), .C(setup_counter_r[0]), .A(n355), .Y(
        n356) );
  NOR2X1 U433 ( .A(setup_counter_r[0]), .B(n353), .Y(N333) );
  NOR2X1 U434 ( .A(n295), .B(n291), .Y(N688) );
  XNOR2XL U435 ( .A(clk_count2[3]), .B(n296), .Y(n295) );
  NOR2X1 U436 ( .A(n106), .B(n293), .Y(n296) );
  NOR2X1 U437 ( .A(n298), .B(n291), .Y(N686) );
  XNOR2XL U438 ( .A(clk_count2[1]), .B(clk_count2[0]), .Y(n298) );
  NOR2X1 U439 ( .A(n290), .B(n291), .Y(N690) );
  AOI22AXL U440 ( .A(i2ccon_o[7]), .B(n292), .D(n293), .C(n294), .Y(n290) );
  OAI21BBX1 U441 ( .A(i2ccon_o[0]), .B(clk_count2[0]), .C(n47), .Y(n292) );
  OAI21BBX1 U442 ( .A(clk_count2[2]), .B(clk_count2[3]), .C(i2ccon_o[7]), .Y(
        n294) );
  AOI211X1 U443 ( .C(n82), .D(n197), .A(n198), .B(n89), .Y(n501) );
  OAI211X1 U444 ( .C(n199), .D(n83), .A(n56), .B(n22), .Y(n198) );
  NAND4X1 U445 ( .A(n200), .B(adrcompen), .C(i2ccon_o[2]), .D(n201), .Y(n197)
         );
  AOI221XL U446 ( .A(n63), .B(fsmsta[4]), .C(n73), .D(n76), .E(n67), .Y(n199)
         );
  NAND4X1 U447 ( .A(n212), .B(n213), .C(n214), .D(n215), .Y(n207) );
  XNOR2XL U448 ( .A(i2cdat_o[3]), .B(i2cadr_o[4]), .Y(n213) );
  XNOR2XL U449 ( .A(i2cdat_o[2]), .B(i2cadr_o[3]), .Y(n212) );
  XNOR2XL U450 ( .A(i2cdat_o[5]), .B(i2cadr_o[6]), .Y(n214) );
  INVX1 U451 ( .A(n254), .Y(n59) );
  AOI32X1 U452 ( .A(n61), .B(n20), .C(n255), .D(n60), .E(sclscl), .Y(n254) );
  INVX1 U453 ( .A(n255), .Y(n60) );
  NAND3X1 U454 ( .A(n87), .B(n20), .C(n61), .Y(n255) );
  INVX1 U455 ( .A(i2ccon_o[3]), .Y(n83) );
  NAND31X1 U456 ( .C(clk_count1[2]), .A(n104), .B(n102), .Y(n308) );
  NAND21X1 U457 ( .B(clkint_ff), .A(clkint), .Y(n280) );
  AOI21X1 U458 ( .B(n86), .C(i2ccon_o[3]), .A(n334), .Y(n327) );
  INVX1 U459 ( .A(sclint), .Y(n86) );
  NAND2X1 U460 ( .A(clkint_ff), .B(n108), .Y(n388) );
  INVX1 U461 ( .A(fsmsync[1]), .Y(n120) );
  NAND2X1 U462 ( .A(bclkcnt[1]), .B(n318), .Y(n313) );
  XOR2X1 U463 ( .A(bclksel), .B(bclkcnt[0]), .Y(n318) );
  NAND3X1 U464 ( .A(fsmsync[0]), .B(n120), .C(fsmsync[2]), .Y(n285) );
  AOI21X1 U465 ( .B(i2ccon_o[0]), .C(i2ccon_o[1]), .A(n41), .Y(n250) );
  INVX1 U466 ( .A(i2ccon_o[6]), .Y(n45) );
  INVX1 U467 ( .A(pedetect), .Y(n87) );
  AND2X1 U468 ( .A(n378), .B(starto_en), .Y(n376) );
  OAI33XL U469 ( .A(n180), .B(n181), .C(n124), .D(n182), .E(n28), .F(n183), 
        .Y(n496) );
  INVX1 U470 ( .A(adrcompen), .Y(n124) );
  OAI21X1 U471 ( .B(n88), .C(n184), .A(n56), .Y(n180) );
  NAND3X1 U472 ( .A(i2ccon_o[0]), .B(n41), .C(i2ccon_o[1]), .Y(n242) );
  INVX1 U473 ( .A(i2ccon_o[4]), .Y(n109) );
  NOR2X1 U474 ( .A(fsmsync[2]), .B(fsmsync[0]), .Y(n289) );
  NOR3XL U475 ( .A(fsmmod[1]), .B(fsmmod[2]), .C(fsmmod[0]), .Y(n228) );
  AOI21X1 U476 ( .B(n286), .C(n287), .A(n267), .Y(N746) );
  AOI211X1 U477 ( .C(n268), .D(n272), .A(n278), .B(n288), .Y(n287) );
  AOI222XL U478 ( .A(n119), .B(n109), .C(i2ccon_o[3]), .D(n273), .E(n118), .F(
        n86), .Y(n286) );
  AOI21AX1 U479 ( .B(sdaint), .C(n117), .A(n270), .Y(n288) );
  AOI21AX1 U480 ( .B(clk_count1[3]), .C(n302), .A(n309), .Y(n240) );
  INVX1 U481 ( .A(clkint), .Y(n108) );
  NOR2X1 U482 ( .A(n113), .B(i2ccon_o[3]), .Y(n375) );
  INVX1 U483 ( .A(clk_count1[0]), .Y(n102) );
  INVX1 U484 ( .A(clk_count1[1]), .Y(n104) );
  AOI32X1 U485 ( .A(n37), .B(i2ccon_o[7]), .C(n248), .D(n249), .E(n250), .Y(
        n247) );
  NOR3XL U486 ( .A(n47), .B(n251), .C(n48), .Y(n248) );
  NAND2X1 U487 ( .A(n289), .B(fsmsync[1]), .Y(n283) );
  NAND3X1 U488 ( .A(nedetect), .B(n113), .C(n327), .Y(n328) );
  INVX1 U489 ( .A(i2ccon_o[7]), .Y(n41) );
  OAI21X1 U490 ( .B(n256), .C(n52), .A(n257), .Y(n507) );
  NOR3XL U491 ( .A(sdai_ff_reg0[0]), .B(sdai_ff_reg0[2]), .C(sdai_ff_reg0[1]), 
        .Y(n256) );
  AOI31X1 U492 ( .A(sdai_ff_reg0[1]), .B(sdai_ff_reg0[0]), .C(sdai_ff_reg0[2]), 
        .D(n28), .Y(n257) );
  OAI21X1 U493 ( .B(n324), .C(n84), .A(n91), .Y(N493) );
  XNOR2XL U494 ( .A(framesync[1]), .B(framesync[0]), .Y(n324) );
  INVX1 U495 ( .A(framesync[2]), .Y(n114) );
  NAND3X1 U496 ( .A(n48), .B(n41), .C(i2ccon_o[1]), .Y(n241) );
  NAND3X1 U497 ( .A(n47), .B(n41), .C(i2ccon_o[0]), .Y(n244) );
  NOR4XL U498 ( .A(n279), .B(n86), .C(n280), .D(n281), .Y(n277) );
  AOI221XL U499 ( .A(fsmmod[0]), .B(n100), .C(n58), .D(n62), .E(n282), .Y(n279) );
  NAND4X1 U500 ( .A(i2ccon_o[6]), .B(n387), .C(n92), .D(n19), .Y(n373) );
  NAND3X1 U501 ( .A(n7), .B(pedetect), .C(n67), .Y(n387) );
  NAND4X1 U502 ( .A(scli_ff_reg0[1]), .B(scli_ff_reg0[0]), .C(n191), .D(n49), 
        .Y(n187) );
  NOR21XL U503 ( .B(scli_ff_reg0[2]), .A(n28), .Y(n191) );
  AOI21X1 U504 ( .B(fsmsta[2]), .C(n66), .A(n79), .Y(n332) );
  INVX1 U505 ( .A(i2ccon_o[1]), .Y(n47) );
  NOR3XL U506 ( .A(n382), .B(i2ccon_o[4]), .C(n388), .Y(n389) );
  INVX1 U507 ( .A(i2ccon_o[0]), .Y(n48) );
  NAND2X1 U508 ( .A(clk_count1[3]), .B(clk_count1[2]), .Y(n309) );
  NOR3XL U509 ( .A(n141), .B(n115), .C(n86), .Y(n490) );
  OAI211X1 U510 ( .C(n107), .D(starto_en), .A(n142), .B(n22), .Y(n141) );
  AOI21X1 U511 ( .B(n265), .C(n266), .A(n267), .Y(N748) );
  AOI221XL U512 ( .A(n110), .B(n268), .C(n269), .D(n86), .E(n270), .Y(n266) );
  AOI22X1 U513 ( .A(i2ccon_o[3]), .B(n273), .C(n119), .D(i2ccon_o[4]), .Y(n265) );
  INVX1 U514 ( .A(n272), .Y(n110) );
  NAND3X1 U515 ( .A(n20), .B(n86), .C(write_data_r), .Y(n354) );
  NOR2X1 U516 ( .A(n308), .B(clk_count1[3]), .Y(n251) );
  OAI211X1 U517 ( .C(fsmsta[0]), .D(n78), .A(n342), .B(n338), .Y(N406) );
  OAI211X1 U518 ( .C(n258), .D(n259), .A(n21), .B(i2ccon_o[6]), .Y(N749) );
  AOI21X1 U519 ( .B(n117), .C(n120), .A(n260), .Y(n259) );
  AOI211X1 U520 ( .C(n78), .D(fsmsta[1]), .A(n261), .B(n83), .Y(n258) );
  OAI211X1 U521 ( .C(fsmsta[4]), .D(n262), .A(n263), .B(n86), .Y(n261) );
  AOI21BX1 U522 ( .C(n396), .B(n397), .A(n188), .Y(N1063) );
  NAND2X1 U523 ( .A(n394), .B(n52), .Y(n397) );
  OAI32X1 U524 ( .A(n394), .B(fsmdet[0]), .C(n52), .D(n395), .E(fsmdet[2]), 
        .Y(n396) );
  AOI31X1 U525 ( .A(n274), .B(n275), .C(n276), .D(n267), .Y(N747) );
  NAND21X1 U526 ( .B(n283), .A(n280), .Y(n275) );
  AOI32X1 U527 ( .A(n120), .B(n121), .C(fsmsync[0]), .D(n284), .E(n83), .Y(
        n274) );
  NOR3XL U528 ( .A(n277), .B(n278), .C(n270), .Y(n276) );
  AOI31X1 U529 ( .A(n379), .B(n380), .C(n381), .D(n373), .Y(N1125) );
  NAND2X1 U530 ( .A(n383), .B(nedetect), .Y(n379) );
  OAI21BBX1 U531 ( .A(i2ccon_o[4]), .B(n375), .C(n57), .Y(n380) );
  AOI31X1 U532 ( .A(n370), .B(n371), .C(n372), .D(n373), .Y(N1126) );
  NAND3X1 U533 ( .A(n57), .B(i2ccon_o[4]), .C(n375), .Y(n371) );
  AOI222XL U534 ( .A(n61), .B(n374), .C(n282), .D(n88), .E(n232), .F(n253), 
        .Y(n372) );
  AOI33X1 U535 ( .A(i2ccon_o[5]), .B(n52), .C(n376), .D(sclint), .E(n377), .F(
        n229), .Y(n370) );
  AOI31X1 U536 ( .A(n384), .B(n385), .C(n386), .D(n373), .Y(N1124) );
  OAI21BBX1 U537 ( .A(n377), .B(sclint), .C(n229), .Y(n385) );
  AOI22X1 U538 ( .A(n383), .B(n88), .C(n61), .D(n374), .Y(n386) );
  AOI33X1 U539 ( .A(n333), .B(n375), .C(n389), .D(n378), .E(i2ccon_o[5]), .F(
        starto_en), .Y(n384) );
  INVX1 U540 ( .A(i2cdat_o[0]), .Y(n81) );
  INVX1 U541 ( .A(i2cdat_o[2]), .Y(n97) );
  INVX1 U542 ( .A(i2cdat_o[1]), .Y(n96) );
  NOR2X1 U543 ( .A(n337), .B(n336), .Y(N470) );
  XNOR2XL U544 ( .A(indelay[1]), .B(indelay[0]), .Y(n337) );
  NOR2X1 U545 ( .A(n316), .B(n317), .Y(N511) );
  XNOR2XL U546 ( .A(bclkcnt[1]), .B(bclkcnt[0]), .Y(n316) );
  NOR2X1 U547 ( .A(bclkcnt[0]), .B(n317), .Y(N510) );
  NOR2X1 U548 ( .A(n392), .B(n188), .Y(N1064) );
  AOI221XL U549 ( .A(fsmdet[2]), .B(fsmdet[0]), .C(n393), .D(n52), .E(n394), 
        .Y(n392) );
  OAI21X1 U550 ( .B(fsmdet[2]), .C(fsmdet[0]), .A(n395), .Y(n393) );
  NOR2X1 U551 ( .A(n391), .B(n188), .Y(N1065) );
  AOI221XL U552 ( .A(sdaint), .B(fsmdet[1]), .C(fsmdet[2]), .D(n94), .E(n90), 
        .Y(n391) );
  NAND4X1 U553 ( .A(n338), .B(n339), .C(n340), .D(n341), .Y(N410) );
  NAND21X1 U554 ( .B(n342), .A(fsmsta[4]), .Y(n339) );
  NAND2X1 U555 ( .A(clk_count1[3]), .B(n308), .Y(n243) );
  INVX1 U556 ( .A(busfree), .Y(n115) );
  INVX1 U557 ( .A(bsd7_tmp), .Y(n98) );
  NOR32XL U558 ( .B(indelay[1]), .C(indelay[2]), .A(indelay[0]), .Y(n271) );
  OAI31XL U559 ( .A(scli_ff_reg0[0]), .B(scli_ff_reg0[2]), .C(scli_ff_reg0[1]), 
        .D(n85), .Y(n190) );
  NAND2X1 U560 ( .A(n178), .B(i2ccon_o[4]), .Y(n272) );
  INVX1 U561 ( .A(nedetect), .Y(n88) );
  INVX1 U562 ( .A(fsmsync[0]), .Y(n117) );
  INVX1 U563 ( .A(fsmsync[2]), .Y(n121) );
  NAND2X1 U564 ( .A(clk_count2[1]), .B(clk_count2[0]), .Y(n293) );
  INVX1 U565 ( .A(adrcomp), .Y(n82) );
  NOR2X1 U566 ( .A(setup_counter_r[1]), .B(setup_counter_r[0]), .Y(n355) );
  ENOX1 U567 ( .A(fsmsync[0]), .B(n121), .C(n271), .D(n260), .Y(n269) );
  INVX1 U568 ( .A(clk_count2[2]), .Y(n106) );
  NAND2X1 U569 ( .A(n107), .B(sclint), .Y(n253) );
  NAND2X1 U570 ( .A(sclscl), .B(pedetect), .Y(n374) );
  OR2X1 U571 ( .A(sdai_ff_reg0[1]), .B(n27), .Y(N433) );
  OR2X1 U572 ( .A(sdai_ff_reg0[0]), .B(n27), .Y(N432) );
  OR2X1 U573 ( .A(sdai_ff), .B(n27), .Y(N431) );
  OR2X1 U574 ( .A(scli_ff), .B(n27), .Y(N412) );
  INVX1 U575 ( .A(clk_count1_ov), .Y(n105) );
  INVX1 U576 ( .A(setup_counter_r[2]), .Y(n99) );
  BUFX3 U577 ( .A(i2ccon_o[3]), .Y(si) );
endmodule


module SNPS_CLOCK_GATE_HIGH_i2c_a0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_i2c_a0_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_i2c_a0_3 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_i2c_a0_4 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_i2c_a0_5 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_i2c_a0_6 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_i2c_a0_7 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_i2c_a0_8 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_i2c_a0_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module extint_a0 ( clkper, rst, newinstr, int0ff, int0ack, int1ff, int1ack, 
        int2ff, iex2ack, int3ff, iex3ack, int4ff, iex4ack, int5ff, iex5ack, 
        int6ff, iex6ack, int7ff, iex7ack, int8ff, iex8ack, int9ff, iex9ack, 
        ie0, it0, ie1, it1, i2fr, iex2, i3fr, iex3, iex4, iex5, iex6, iex7, 
        iex8, iex9, iex10, iex11, iex12, sfraddr, sfrdatai, sfrwe );
  input [6:0] sfraddr;
  input [7:0] sfrdatai;
  input clkper, rst, newinstr, int0ff, int0ack, int1ff, int1ack, int2ff,
         iex2ack, int3ff, iex3ack, int4ff, iex4ack, int5ff, iex5ack, int6ff,
         iex6ack, int7ff, iex7ack, int8ff, iex8ack, int9ff, iex9ack, sfrwe;
  output ie0, it0, ie1, it1, i2fr, iex2, i3fr, iex3, iex4, iex5, iex6, iex7,
         iex8, iex9, iex10, iex11, iex12;
  wire   int0_ff1, int0_fall, int0_clr, N23, int1_ff1, int1_fall, int1_clr,
         N51, int2_ff1, iex2_set, N71, int3_ff1, iex3_set, N90, iex4_set,
         int4_ff1, iex5_set, int5_ff1, iex6_set, int6_ff1, iex7_set, int7_ff1,
         iex8_set, int8_ff1, iex9_set, int9_ff1, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129;

  DFFQX1 int4_ff1_reg ( .D(n24), .C(clkper), .Q(int4_ff1) );
  DFFQX1 int5_ff1_reg ( .D(n16), .C(clkper), .Q(int5_ff1) );
  DFFQX1 int6_ff1_reg ( .D(n22), .C(clkper), .Q(int6_ff1) );
  DFFQX1 int7_ff1_reg ( .D(n23), .C(clkper), .Q(int7_ff1) );
  DFFQX1 int8_ff1_reg ( .D(n127), .C(clkper), .Q(int8_ff1) );
  DFFQX1 int9_ff1_reg ( .D(n14), .C(clkper), .Q(int9_ff1) );
  DFFQX1 iex2_set_reg ( .D(n110), .C(clkper), .Q(iex2_set) );
  DFFQX1 iex3_set_reg ( .D(n107), .C(clkper), .Q(iex3_set) );
  DFFQX1 iex4_set_reg ( .D(n105), .C(clkper), .Q(iex4_set) );
  DFFQX1 iex5_set_reg ( .D(n103), .C(clkper), .Q(iex5_set) );
  DFFQX1 iex6_set_reg ( .D(n101), .C(clkper), .Q(iex6_set) );
  DFFQX1 iex7_set_reg ( .D(n99), .C(clkper), .Q(iex7_set) );
  DFFQX1 iex8_set_reg ( .D(n97), .C(clkper), .Q(iex8_set) );
  DFFQX1 iex9_set_reg ( .D(n95), .C(clkper), .Q(iex9_set) );
  DFFQX1 int0_fall_reg ( .D(n116), .C(clkper), .Q(int0_fall) );
  DFFQX1 int1_fall_reg ( .D(n112), .C(clkper), .Q(int1_fall) );
  DFFQX1 int2_ff1_reg ( .D(N71), .C(clkper), .Q(int2_ff1) );
  DFFQX1 int3_ff1_reg ( .D(N90), .C(clkper), .Q(int3_ff1) );
  DFFQX1 int0_clr_reg ( .D(n118), .C(clkper), .Q(int0_clr) );
  DFFQX1 int1_clr_reg ( .D(n114), .C(clkper), .Q(int1_clr) );
  DFFQX1 int0_ff1_reg ( .D(N23), .C(clkper), .Q(int0_ff1) );
  DFFQX1 int1_ff1_reg ( .D(N51), .C(clkper), .Q(int1_ff1) );
  DFFQX1 iex8_s_reg ( .D(n96), .C(clkper), .Q(iex8) );
  DFFQX1 iex9_s_reg ( .D(n94), .C(clkper), .Q(iex9) );
  DFFQX1 iex5_s_reg ( .D(n102), .C(clkper), .Q(iex5) );
  DFFQX1 iex6_s_reg ( .D(n100), .C(clkper), .Q(iex6) );
  DFFQX1 iex4_s_reg ( .D(n104), .C(clkper), .Q(iex4) );
  DFFQX1 iex2_s_reg ( .D(n109), .C(clkper), .Q(iex2) );
  DFFQX1 iex7_s_reg ( .D(n98), .C(clkper), .Q(iex7) );
  DFFQX1 ie0_s_reg ( .D(n115), .C(clkper), .Q(ie0) );
  DFFQX1 ie1_s_reg ( .D(n111), .C(clkper), .Q(ie1) );
  DFFQX1 iex3_s_reg ( .D(n106), .C(clkper), .Q(iex3) );
  DFFQX1 it1_s_reg ( .D(n113), .C(clkper), .Q(it1) );
  DFFQX1 i2fr_s_reg ( .D(n18), .C(clkper), .Q(i2fr) );
  DFFQX1 it0_s_reg ( .D(n117), .C(clkper), .Q(it0) );
  DFFQX1 i3fr_s_reg ( .D(n108), .C(clkper), .Q(i3fr) );
  INVX1 U3 ( .A(1'b1), .Y(iex12) );
  INVX1 U5 ( .A(1'b1), .Y(iex11) );
  INVX1 U7 ( .A(1'b1), .Y(iex10) );
  NOR2X1 U9 ( .A(newinstr), .B(rst), .Y(n47) );
  INVX1 U10 ( .A(n47), .Y(n7) );
  INVX1 U11 ( .A(n47), .Y(n8) );
  NOR2X1 U12 ( .A(n10), .B(n20), .Y(n56) );
  INVX1 U13 ( .A(n57), .Y(n20) );
  INVX1 U14 ( .A(n81), .Y(n17) );
  INVX1 U15 ( .A(n77), .Y(n19) );
  INVX1 U16 ( .A(n46), .Y(n21) );
  INVX1 U17 ( .A(n12), .Y(n10) );
  INVX1 U18 ( .A(n13), .Y(n11) );
  NAND32X1 U19 ( .B(sfraddr[3]), .C(n9), .A(n74), .Y(n57) );
  AOI31X1 U20 ( .A(sfraddr[6]), .B(sfraddr[3]), .C(n74), .D(n10), .Y(n77) );
  NOR42XL U21 ( .C(sfrwe), .D(n93), .A(sfraddr[0]), .B(sfraddr[1]), .Y(n74) );
  NOR3XL U22 ( .A(sfraddr[2]), .B(sfraddr[5]), .C(sfraddr[4]), .Y(n93) );
  NAND2X1 U23 ( .A(n51), .B(n52), .Y(n46) );
  NOR43XL U24 ( .B(sfraddr[2]), .C(sfraddr[0]), .D(sfraddr[1]), .A(sfraddr[6]), 
        .Y(n52) );
  AND4X1 U25 ( .A(sfraddr[3]), .B(sfraddr[4]), .C(sfraddr[5]), .D(sfrwe), .Y(
        n51) );
  NAND3X1 U26 ( .A(sfraddr[3]), .B(n9), .C(n74), .Y(n81) );
  INVX1 U27 ( .A(sfraddr[6]), .Y(n9) );
  INVX1 U28 ( .A(n58), .Y(n23) );
  NAND2X1 U29 ( .A(n13), .B(n15), .Y(N71) );
  INVX1 U30 ( .A(int0ack), .Y(n42) );
  INVX1 U31 ( .A(int1ack), .Y(n43) );
  INVX1 U32 ( .A(rst), .Y(n12) );
  NAND2X1 U33 ( .A(n13), .B(n25), .Y(N90) );
  INVX1 U34 ( .A(n53), .Y(n127) );
  INVX1 U35 ( .A(n64), .Y(n16) );
  OAI21X1 U36 ( .B(n34), .C(n19), .A(n71), .Y(n108) );
  NAND3X1 U37 ( .A(n19), .B(n13), .C(sfrdatai[6]), .Y(n71) );
  INVX1 U38 ( .A(n67), .Y(n24) );
  INVX1 U39 ( .A(n48), .Y(n14) );
  OAI32X1 U40 ( .A(n27), .B(int0ack), .C(n7), .D(n10), .E(n91), .Y(n116) );
  OAI32X1 U41 ( .A(n29), .B(int1ack), .C(n7), .D(n10), .E(n84), .Y(n112) );
  OAI22X1 U42 ( .A(n11), .B(n43), .C(n8), .D(n28), .Y(n114) );
  OAI22X1 U43 ( .A(n11), .B(n42), .C(n8), .D(n26), .Y(n118) );
  NAND2X1 U44 ( .A(int7ff), .B(n13), .Y(n58) );
  INVX1 U45 ( .A(int2ff), .Y(n15) );
  INVX1 U46 ( .A(int3ff), .Y(n25) );
  INVX1 U47 ( .A(n61), .Y(n22) );
  NAND2X1 U48 ( .A(int8ff), .B(n12), .Y(n53) );
  NOR2X1 U49 ( .A(n10), .B(n129), .Y(N51) );
  NOR2X1 U50 ( .A(n10), .B(n128), .Y(N23) );
  NAND2X1 U51 ( .A(int5ff), .B(n12), .Y(n64) );
  OAI32X1 U52 ( .A(n37), .B(iex5ack), .C(n7), .D(int5_ff1), .E(n64), .Y(n103)
         );
  INVX1 U53 ( .A(iex5_set), .Y(n37) );
  GEN2XL U54 ( .D(n17), .E(sfrdatai[3]), .C(n78), .B(n13), .A(n79), .Y(n111)
         );
  NOR4XL U55 ( .A(n80), .B(int1_clr), .C(n10), .D(int1ack), .Y(n79) );
  OAI31XL U56 ( .A(n17), .B(it1), .C(int1ff), .D(n82), .Y(n78) );
  NAND3X1 U57 ( .A(it1), .B(n81), .C(ie1), .Y(n80) );
  GEN2XL U58 ( .D(n17), .E(sfrdatai[1]), .C(n86), .B(n13), .A(n87), .Y(n115)
         );
  NOR4XL U59 ( .A(n88), .B(int0_clr), .C(n10), .D(int0ack), .Y(n87) );
  OAI31XL U60 ( .A(n17), .B(it0), .C(int0ff), .D(n89), .Y(n86) );
  NAND3X1 U61 ( .A(it0), .B(n81), .C(ie0), .Y(n88) );
  NAND2X1 U62 ( .A(int4ff), .B(n12), .Y(n67) );
  OAI32X1 U63 ( .A(n36), .B(iex4ack), .C(n7), .D(int4_ff1), .E(n67), .Y(n105)
         );
  INVX1 U64 ( .A(iex4_set), .Y(n36) );
  NOR2X1 U65 ( .A(n10), .B(n92), .Y(n117) );
  AOI22X1 U66 ( .A(it0), .B(n81), .C(n17), .D(sfrdatai[0]), .Y(n92) );
  NOR2X1 U67 ( .A(n10), .B(n85), .Y(n113) );
  AOI22X1 U68 ( .A(it1), .B(n81), .C(n17), .D(sfrdatai[2]), .Y(n85) );
  OAI21X1 U69 ( .B(n11), .C(n44), .A(n45), .Y(n94) );
  NAND4X1 U70 ( .A(iex9), .B(n46), .C(n125), .D(n12), .Y(n45) );
  AOI32X1 U71 ( .A(n46), .B(n125), .C(iex9_set), .D(sfrdatai[1]), .E(n21), .Y(
        n44) );
  INVX1 U72 ( .A(iex9ack), .Y(n125) );
  OAI21X1 U73 ( .B(rst), .C(n49), .A(n50), .Y(n96) );
  NAND4X1 U74 ( .A(iex8), .B(n46), .C(n126), .D(n13), .Y(n50) );
  AOI32X1 U75 ( .A(n46), .B(n126), .C(iex8_set), .D(sfrdatai[0]), .E(n21), .Y(
        n49) );
  INVX1 U76 ( .A(iex8ack), .Y(n126) );
  OAI21X1 U77 ( .B(rst), .C(n54), .A(n55), .Y(n98) );
  NAND3X1 U78 ( .A(n56), .B(n119), .C(iex7), .Y(n55) );
  AOI32X1 U79 ( .A(n57), .B(n119), .C(iex7_set), .D(n20), .E(sfrdatai[0]), .Y(
        n54) );
  INVX1 U80 ( .A(iex7ack), .Y(n119) );
  OAI21X1 U81 ( .B(n11), .C(n59), .A(n60), .Y(n100) );
  NAND3X1 U82 ( .A(n56), .B(n124), .C(iex6), .Y(n60) );
  AOI32X1 U83 ( .A(n57), .B(n124), .C(iex6_set), .D(sfrdatai[5]), .E(n20), .Y(
        n59) );
  INVX1 U84 ( .A(iex6ack), .Y(n124) );
  OAI21X1 U85 ( .B(n11), .C(n62), .A(n63), .Y(n102) );
  NAND3X1 U86 ( .A(n56), .B(n123), .C(iex5), .Y(n63) );
  AOI32X1 U87 ( .A(n57), .B(n123), .C(iex5_set), .D(sfrdatai[4]), .E(n20), .Y(
        n62) );
  INVX1 U88 ( .A(iex5ack), .Y(n123) );
  OAI21X1 U89 ( .B(n11), .C(n65), .A(n66), .Y(n104) );
  NAND3X1 U90 ( .A(n56), .B(n122), .C(iex4), .Y(n66) );
  AOI32X1 U91 ( .A(n57), .B(n122), .C(iex4_set), .D(sfrdatai[3]), .E(n20), .Y(
        n65) );
  INVX1 U92 ( .A(iex4ack), .Y(n122) );
  OAI21X1 U93 ( .B(n11), .C(n68), .A(n69), .Y(n106) );
  NAND3X1 U94 ( .A(n56), .B(n121), .C(iex3), .Y(n69) );
  AOI32X1 U95 ( .A(n57), .B(n121), .C(iex3_set), .D(sfrdatai[2]), .E(n20), .Y(
        n68) );
  INVX1 U96 ( .A(iex3ack), .Y(n121) );
  OAI21X1 U97 ( .B(n11), .C(n72), .A(n73), .Y(n109) );
  NAND3X1 U98 ( .A(n56), .B(n120), .C(iex2), .Y(n73) );
  AOI32X1 U99 ( .A(n57), .B(n120), .C(iex2_set), .D(n20), .E(sfrdatai[1]), .Y(
        n72) );
  INVX1 U100 ( .A(iex2ack), .Y(n120) );
  NAND4X1 U101 ( .A(n28), .B(n43), .C(n81), .D(n83), .Y(n82) );
  AOI21AX1 U102 ( .B(n29), .C(n84), .A(it1), .Y(n83) );
  NAND4X1 U103 ( .A(n26), .B(n42), .C(n81), .D(n90), .Y(n89) );
  AOI21AX1 U104 ( .B(n27), .C(n91), .A(it0), .Y(n90) );
  INVX1 U105 ( .A(n76), .Y(n18) );
  AOI32X1 U106 ( .A(sfrdatai[5]), .B(n12), .C(n19), .D(n77), .E(i2fr), .Y(n76)
         );
  NAND2X1 U107 ( .A(int9ff), .B(n13), .Y(n48) );
  INVX1 U108 ( .A(rst), .Y(n13) );
  OAI32X1 U109 ( .A(n8), .B(iex9ack), .C(n41), .D(int9_ff1), .E(n48), .Y(n95)
         );
  INVX1 U110 ( .A(iex9_set), .Y(n41) );
  OAI32X1 U111 ( .A(n39), .B(iex7ack), .C(n7), .D(int7_ff1), .E(n58), .Y(n99)
         );
  INVX1 U112 ( .A(iex7_set), .Y(n39) );
  OAI32X1 U113 ( .A(n40), .B(iex8ack), .C(n7), .D(int8_ff1), .E(n53), .Y(n97)
         );
  INVX1 U114 ( .A(iex8_set), .Y(n40) );
  OAI32X1 U115 ( .A(n38), .B(iex6ack), .C(n8), .D(int6_ff1), .E(n61), .Y(n101)
         );
  INVX1 U116 ( .A(iex6_set), .Y(n38) );
  OAI32X1 U117 ( .A(n35), .B(iex3ack), .C(n8), .D(n11), .E(n70), .Y(n107) );
  INVX1 U118 ( .A(iex3_set), .Y(n35) );
  AOI33X1 U119 ( .A(n34), .B(n25), .C(int3_ff1), .D(i3fr), .E(n33), .F(int3ff), 
        .Y(n70) );
  INVX1 U120 ( .A(int3_ff1), .Y(n33) );
  OAI32X1 U121 ( .A(n32), .B(iex2ack), .C(n8), .D(n11), .E(n75), .Y(n110) );
  INVX1 U122 ( .A(iex2_set), .Y(n32) );
  AOI33X1 U123 ( .A(n31), .B(n15), .C(int2_ff1), .D(i2fr), .E(n30), .F(int2ff), 
        .Y(n75) );
  INVX1 U124 ( .A(int2_ff1), .Y(n30) );
  NAND2X1 U125 ( .A(int6ff), .B(n13), .Y(n61) );
  INVX1 U126 ( .A(int0ff), .Y(n128) );
  INVX1 U127 ( .A(int1ff), .Y(n129) );
  NAND2X1 U128 ( .A(int1_ff1), .B(n129), .Y(n84) );
  NAND2X1 U129 ( .A(int0_ff1), .B(n128), .Y(n91) );
  INVX1 U130 ( .A(int1_clr), .Y(n28) );
  INVX1 U131 ( .A(int0_clr), .Y(n26) );
  INVX1 U132 ( .A(i3fr), .Y(n34) );
  INVX1 U133 ( .A(i2fr), .Y(n31) );
  INVX1 U134 ( .A(int1_fall), .Y(n29) );
  INVX1 U135 ( .A(int0_fall), .Y(n27) );
endmodule


module isr_a0 ( clkper, rst, intcall, retiinstr, int_vect_03, int_vect_0b, 
        t0ff, int_vect_13, int_vect_1b, t1ff, int_vect_23, i2c_int, rxd0ff, 
        int_vect_43, sdaiff, int_vect_4b, int_vect_53, int_vect_5b, 
        int_vect_63, int_vect_6b, int_vect_8b, int_vect_93, int_vect_9b, 
        int_vect_a3, int_vect_ab, irq, intvect, int_ack_03, int_ack_0b, 
        int_ack_13, int_ack_1b, int_ack_43, int_ack_4b, int_ack_53, int_ack_5b, 
        int_ack_63, int_ack_6b, int_ack_8b, int_ack_93, int_ack_9b, int_ack_a3, 
        int_ack_ab, is_reg, ip0, ip1, ien0, ien1, ien2, isr_tm, sfraddr, 
        sfrdatai, sfrwe );
  output [4:0] intvect;
  output [3:0] is_reg;
  output [5:0] ip0;
  output [5:0] ip1;
  output [7:0] ien0;
  output [5:0] ien1;
  output [5:0] ien2;
  input [6:0] sfraddr;
  input [7:0] sfrdatai;
  input clkper, rst, intcall, retiinstr, int_vect_03, int_vect_0b, t0ff,
         int_vect_13, int_vect_1b, t1ff, int_vect_23, i2c_int, rxd0ff,
         int_vect_43, sdaiff, int_vect_4b, int_vect_53, int_vect_5b,
         int_vect_63, int_vect_6b, int_vect_8b, int_vect_93, int_vect_9b,
         int_vect_a3, int_vect_ab, sfrwe;
  output irq, int_ack_03, int_ack_0b, int_ack_13, int_ack_1b, int_ack_43,
         int_ack_4b, int_ack_53, int_ack_5b, int_ack_63, int_ack_6b,
         int_ack_8b, int_ack_93, int_ack_9b, int_ack_a3, int_ack_ab, isr_tm;
  wire   N38, N39, N40, N41, N42, N43, N44, N45, N49, N50, N51, N52, N53, N54,
         N55, N58, N59, N60, N61, N62, N63, N64, N67, N68, N69, N70, N71, N72,
         N73, N76, N77, N78, N79, N80, N81, N82, irq_r, N200, N207, N208, N209,
         N210, N211, N212, net12106, net12112, net12117, net12122, net12127,
         net12132, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n201, n202, n203;

  SNPS_CLOCK_GATE_HIGH_isr_a0_0 clk_gate_ien0_reg_reg ( .CLK(clkper), .EN(N38), 
        .ENCLK(net12106), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_isr_a0_5 clk_gate_ien1_reg_reg ( .CLK(clkper), .EN(N49), 
        .ENCLK(net12112), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_isr_a0_4 clk_gate_ien2_reg_reg ( .CLK(clkper), .EN(N58), 
        .ENCLK(net12117), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_isr_a0_3 clk_gate_ip0_reg_reg ( .CLK(clkper), .EN(N67), 
        .ENCLK(net12122), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_isr_a0_2 clk_gate_ip1_reg_reg ( .CLK(clkper), .EN(N76), 
        .ENCLK(net12127), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_isr_a0_1 clk_gate_intvect_reg_reg ( .CLK(clkper), .EN(
        N207), .ENCLK(net12132), .TE(1'b0) );
  DFFQX1 intvect_reg_reg_4_ ( .D(N212), .C(net12132), .Q(intvect[4]) );
  DFFQX1 intvect_reg_reg_3_ ( .D(N211), .C(net12132), .Q(intvect[3]) );
  DFFQX1 intvect_reg_reg_2_ ( .D(N210), .C(net12132), .Q(intvect[2]) );
  DFFQX1 intvect_reg_reg_1_ ( .D(N209), .C(net12132), .Q(intvect[1]) );
  DFFQX1 intvect_reg_reg_0_ ( .D(N208), .C(net12132), .Q(intvect[0]) );
  DFFQX1 is_reg_s_reg_0_ ( .D(n199), .C(clkper), .Q(is_reg[0]) );
  DFFQX1 is_reg_s_reg_1_ ( .D(n196), .C(clkper), .Q(is_reg[1]) );
  DFFQX1 is_reg_s_reg_2_ ( .D(n197), .C(clkper), .Q(is_reg[2]) );
  DFFQX1 is_reg_s_reg_3_ ( .D(n198), .C(clkper), .Q(is_reg[3]) );
  DFFQX1 irq_r_reg ( .D(N200), .C(clkper), .Q(irq_r) );
  DFFQX1 ien0_reg_reg_4_ ( .D(N43), .C(net12106), .Q(ien0[4]) );
  DFFQX1 ien0_reg_reg_3_ ( .D(N42), .C(net12106), .Q(ien0[3]) );
  DFFQX1 ien0_reg_reg_1_ ( .D(N40), .C(net12106), .Q(ien0[1]) );
  DFFQX1 ien2_reg_reg_2_ ( .D(N61), .C(net12117), .Q(ien2[2]) );
  DFFQX1 ien0_reg_reg_5_ ( .D(N44), .C(net12106), .Q(ien0[5]) );
  DFFQX1 ien2_reg_reg_3_ ( .D(N62), .C(net12117), .Q(ien2[3]) );
  DFFQX1 ien0_reg_reg_2_ ( .D(N41), .C(net12106), .Q(ien0[2]) );
  DFFQX1 ien2_reg_reg_1_ ( .D(N60), .C(net12117), .Q(ien2[1]) );
  DFFQX1 ien1_reg_reg_2_ ( .D(N52), .C(net12112), .Q(ien1[2]) );
  DFFQX1 ip1_reg_reg_2_ ( .D(N79), .C(net12127), .Q(ip1[2]) );
  DFFQX1 ien2_reg_reg_0_ ( .D(N59), .C(net12117), .Q(ien2[0]) );
  DFFQX1 ien1_reg_reg_0_ ( .D(N50), .C(net12112), .Q(ien1[0]) );
  DFFQX1 ien2_reg_reg_5_ ( .D(N64), .C(net12117), .Q(ien2[5]) );
  DFFQX1 ien1_reg_reg_3_ ( .D(N53), .C(net12112), .Q(ien1[3]) );
  DFFQX1 ien1_reg_reg_4_ ( .D(N54), .C(net12112), .Q(ien1[4]) );
  DFFQX1 ien1_reg_reg_5_ ( .D(N55), .C(net12112), .Q(ien1[5]) );
  DFFQX1 ien1_reg_reg_1_ ( .D(N51), .C(net12112), .Q(ien1[1]) );
  DFFQX1 ien2_reg_reg_4_ ( .D(N63), .C(net12117), .Q(ien2[4]) );
  DFFQX1 ien0_reg_reg_0_ ( .D(N39), .C(net12106), .Q(ien0[0]) );
  DFFQX1 ien0_reg_reg_6_ ( .D(N45), .C(net12106), .Q(ien0[7]) );
  DFFQX1 ip1_reg_reg_1_ ( .D(N78), .C(net12127), .Q(ip1[1]) );
  DFFQX1 ip1_reg_reg_3_ ( .D(N80), .C(net12127), .Q(ip1[3]) );
  DFFQX1 ip1_reg_reg_5_ ( .D(N82), .C(net12127), .Q(ip1[5]) );
  DFFQX1 isr_tm_reg_reg ( .D(n200), .C(clkper), .Q(isr_tm) );
  DFFQX1 ip0_reg_reg_1_ ( .D(N69), .C(net12122), .Q(ip0[1]) );
  DFFQX1 ip0_reg_reg_5_ ( .D(N73), .C(net12122), .Q(ip0[5]) );
  DFFQX1 ip0_reg_reg_3_ ( .D(N71), .C(net12122), .Q(ip0[3]) );
  DFFQX1 ip0_reg_reg_4_ ( .D(N72), .C(net12122), .Q(ip0[4]) );
  DFFQX1 ip1_reg_reg_4_ ( .D(N81), .C(net12127), .Q(ip1[4]) );
  DFFQX1 ip1_reg_reg_0_ ( .D(N77), .C(net12127), .Q(ip1[0]) );
  DFFQX1 ip0_reg_reg_0_ ( .D(N68), .C(net12122), .Q(ip0[0]) );
  DFFQX1 ip0_reg_reg_2_ ( .D(N70), .C(net12122), .Q(ip0[2]) );
  INVX1 U3 ( .A(1'b1), .Y(ien0[6]) );
  NAND3X1 U5 ( .A(n3), .B(n5), .C(n78), .Y(n83) );
  NAND3X1 U6 ( .A(n78), .B(n3), .C(n4), .Y(n82) );
  NAND3X1 U7 ( .A(sfraddr[0]), .B(n5), .C(n78), .Y(n79) );
  NAND3X1 U8 ( .A(n78), .B(sfraddr[0]), .C(n4), .Y(n77) );
  NOR2X1 U9 ( .A(n6), .B(n83), .Y(N39) );
  NOR2X1 U10 ( .A(n7), .B(n83), .Y(N40) );
  NOR2X1 U11 ( .A(n8), .B(n83), .Y(N41) );
  NOR2X1 U12 ( .A(n9), .B(n83), .Y(N42) );
  NOR2X1 U13 ( .A(n10), .B(n83), .Y(N43) );
  NOR2X1 U14 ( .A(n11), .B(n83), .Y(N44) );
  NOR2X1 U15 ( .A(n77), .B(n6), .Y(N77) );
  NOR2X1 U16 ( .A(n77), .B(n7), .Y(N78) );
  NOR2X1 U17 ( .A(n77), .B(n8), .Y(N79) );
  NOR2X1 U18 ( .A(n77), .B(n9), .Y(N80) );
  NOR2X1 U19 ( .A(n77), .B(n10), .Y(N81) );
  NOR2X1 U20 ( .A(n11), .B(n77), .Y(N82) );
  NOR2X1 U21 ( .A(n6), .B(n79), .Y(N68) );
  NOR2X1 U22 ( .A(n7), .B(n79), .Y(N69) );
  NOR2X1 U23 ( .A(n8), .B(n79), .Y(N70) );
  NOR2X1 U24 ( .A(n9), .B(n79), .Y(N71) );
  NOR2X1 U25 ( .A(n10), .B(n79), .Y(N72) );
  NOR2X1 U26 ( .A(n11), .B(n79), .Y(N73) );
  NOR2X1 U27 ( .A(n6), .B(n80), .Y(N59) );
  NOR2X1 U28 ( .A(n7), .B(n80), .Y(N60) );
  NOR2X1 U29 ( .A(n8), .B(n80), .Y(N61) );
  NOR2X1 U30 ( .A(n9), .B(n80), .Y(N62) );
  NOR2X1 U31 ( .A(n10), .B(n80), .Y(N63) );
  NOR2X1 U32 ( .A(n11), .B(n80), .Y(N64) );
  NOR2X1 U33 ( .A(n6), .B(n82), .Y(N50) );
  NOR2X1 U34 ( .A(n7), .B(n82), .Y(N51) );
  NOR2X1 U35 ( .A(n8), .B(n82), .Y(N52) );
  NOR2X1 U36 ( .A(n9), .B(n82), .Y(N53) );
  NOR2X1 U37 ( .A(n10), .B(n82), .Y(N54) );
  NOR2X1 U38 ( .A(n11), .B(n82), .Y(N55) );
  NAND2X1 U39 ( .A(n12), .B(n80), .Y(N58) );
  NAND2X1 U40 ( .A(n12), .B(n77), .Y(N76) );
  NAND2X1 U41 ( .A(n12), .B(n82), .Y(N49) );
  NAND2X1 U42 ( .A(n12), .B(n79), .Y(N67) );
  NAND2X1 U43 ( .A(n12), .B(n83), .Y(N38) );
  INVX1 U44 ( .A(n5), .Y(n4) );
  INVX1 U45 ( .A(sfraddr[0]), .Y(n3) );
  NOR32XL U46 ( .B(n106), .C(n107), .A(n108), .Y(n92) );
  AND4X1 U47 ( .A(n107), .B(n88), .C(n114), .D(n109), .Y(n85) );
  NOR21XL U48 ( .B(n97), .A(n105), .Y(n114) );
  NAND2X1 U49 ( .A(n203), .B(n12), .Y(n43) );
  INVX1 U50 ( .A(n48), .Y(n202) );
  INVX1 U51 ( .A(n121), .Y(n16) );
  NAND31X1 U52 ( .C(sfraddr[6]), .A(n12), .B(sfrwe), .Y(n70) );
  NOR21XL U53 ( .B(sfrdatai[7]), .A(n83), .Y(N45) );
  NAND4X1 U54 ( .A(sfraddr[3]), .B(sfraddr[1]), .C(n4), .D(n81), .Y(n80) );
  NOR4XL U55 ( .A(sfraddr[5]), .B(sfraddr[2]), .C(sfraddr[0]), .D(n70), .Y(n81) );
  AND3X1 U56 ( .A(sfraddr[5]), .B(sfraddr[3]), .C(n84), .Y(n78) );
  NOR3XL U57 ( .A(n70), .B(sfraddr[2]), .C(sfraddr[1]), .Y(n84) );
  INVX1 U58 ( .A(sfraddr[4]), .Y(n5) );
  INVX1 U59 ( .A(sfrdatai[5]), .Y(n11) );
  INVX1 U60 ( .A(sfrdatai[0]), .Y(n6) );
  INVX1 U61 ( .A(sfrdatai[1]), .Y(n7) );
  INVX1 U62 ( .A(sfrdatai[2]), .Y(n8) );
  INVX1 U63 ( .A(sfrdatai[3]), .Y(n9) );
  INVX1 U64 ( .A(sfrdatai[4]), .Y(n10) );
  NOR32XL U65 ( .B(n113), .C(n112), .A(n127), .Y(n125) );
  NOR32XL U66 ( .B(n91), .C(n93), .A(n90), .Y(n117) );
  NOR32XL U67 ( .B(n126), .C(n117), .A(n116), .Y(n119) );
  NAND31X1 U68 ( .C(n124), .A(n129), .B(n125), .Y(n90) );
  NOR43XL U69 ( .B(n98), .C(n123), .D(n106), .A(n104), .Y(n86) );
  AOI21X1 U70 ( .B(n127), .C(n112), .A(n128), .Y(n123) );
  AOI21X1 U71 ( .B(n93), .C(n91), .A(n90), .Y(n128) );
  NOR32XL U72 ( .B(n94), .C(n96), .A(n95), .Y(n112) );
  NOR21XL U73 ( .B(n182), .A(n153), .Y(n175) );
  NOR21XL U74 ( .B(n184), .A(n144), .Y(n159) );
  OAI211X1 U75 ( .C(n90), .D(n93), .A(n109), .B(n110), .Y(n101) );
  NAND21X1 U76 ( .B(n126), .A(n117), .Y(n106) );
  NAND21X1 U77 ( .B(n118), .A(n119), .Y(n97) );
  AND2X1 U78 ( .A(n116), .B(n117), .Y(n105) );
  NAND2X1 U79 ( .A(n119), .B(n118), .Y(n121) );
  NAND2X1 U80 ( .A(n159), .B(n183), .Y(n153) );
  NOR3XL U81 ( .A(n130), .B(rst), .C(intcall), .Y(N200) );
  NOR4XL U82 ( .A(n115), .B(n120), .C(n122), .D(n121), .Y(n130) );
  AOI31X1 U83 ( .A(n97), .B(n98), .C(n99), .D(rst), .Y(N209) );
  NOR2X1 U84 ( .A(n100), .B(n101), .Y(n99) );
  AOI31X1 U85 ( .A(n87), .B(n88), .C(n14), .D(rst), .Y(N210) );
  NAND32X1 U86 ( .B(n94), .C(n95), .A(n96), .Y(n87) );
  INVX1 U87 ( .A(n89), .Y(n14) );
  OAI31XL U88 ( .A(n90), .B(n19), .C(n91), .D(n92), .Y(n89) );
  AOI31X1 U89 ( .A(n15), .B(n92), .C(n102), .D(rst), .Y(N208) );
  INVX1 U90 ( .A(n101), .Y(n15) );
  NOR3XL U91 ( .A(n103), .B(n104), .C(n105), .Y(n102) );
  NOR2X1 U92 ( .A(rst), .B(n86), .Y(N211) );
  NOR2X1 U93 ( .A(rst), .B(n85), .Y(N212) );
  NAND4X1 U94 ( .A(n86), .B(n96), .C(n85), .D(n111), .Y(N207) );
  NOR43XL U95 ( .B(n94), .C(n110), .D(n12), .A(n108), .Y(n111) );
  NAND2X1 U96 ( .A(n175), .B(n176), .Y(n167) );
  NOR21XL U97 ( .B(n112), .A(n113), .Y(n108) );
  NAND21X1 U98 ( .B(n129), .A(n125), .Y(n98) );
  AND2X1 U99 ( .A(n124), .B(n125), .Y(n104) );
  NAND2X1 U100 ( .A(n95), .B(n96), .Y(n110) );
  INVX1 U101 ( .A(n93), .Y(n19) );
  NAND31X1 U102 ( .C(retiinstr), .A(n202), .B(n12), .Y(n47) );
  INVX1 U103 ( .A(intcall), .Y(n203) );
  INVX1 U104 ( .A(rst), .Y(n12) );
  NOR2X1 U105 ( .A(n203), .B(rst), .Y(n48) );
  NAND42X1 U106 ( .C(n120), .D(n121), .A(n122), .B(n18), .Y(n107) );
  NAND3X1 U107 ( .A(n16), .B(n18), .C(n120), .Y(n88) );
  NAND2X1 U108 ( .A(n115), .B(n16), .Y(n109) );
  INVX1 U109 ( .A(n115), .Y(n18) );
  OAI32X1 U110 ( .A(n31), .B(rst), .C(n13), .D(n68), .E(n11), .Y(n200) );
  INVX1 U111 ( .A(n68), .Y(n13) );
  NAND4XL U112 ( .A(sfraddr[1]), .B(sfraddr[0]), .C(sfraddr[2]), .D(n69), .Y(
        n68) );
  NOR4XL U113 ( .A(sfraddr[5]), .B(n4), .C(sfraddr[3]), .D(n70), .Y(n69) );
  NOR21XL U114 ( .B(n192), .A(n161), .Y(n155) );
  NOR21XL U115 ( .B(n190), .A(n187), .Y(n178) );
  AOI211X1 U116 ( .C(n136), .D(n139), .A(n103), .B(n100), .Y(n96) );
  AOI21BBXL U117 ( .B(n182), .C(n24), .A(n151), .Y(n180) );
  AOI21BBXL U118 ( .B(n184), .C(n26), .A(n142), .Y(n157) );
  AOI21BBXL U119 ( .B(n25), .C(n192), .A(n160), .Y(n154) );
  AOI21BBXL U120 ( .B(n23), .C(n190), .A(n186), .Y(n177) );
  OAI222XL U121 ( .A(n20), .B(n17), .C(n166), .D(n167), .E(n168), .F(n27), .Y(
        n149) );
  AOI21BBXL U122 ( .B(n169), .C(n20), .A(n170), .Y(n168) );
  INVX1 U123 ( .A(n171), .Y(n17) );
  AND2X1 U124 ( .A(n178), .B(n189), .Y(n170) );
  AND3X1 U125 ( .A(n133), .B(n141), .C(n156), .Y(n183) );
  OAI21X1 U126 ( .B(n24), .C(n191), .A(n154), .Y(n186) );
  OAI21X1 U127 ( .B(n183), .C(n25), .A(n157), .Y(n151) );
  OAI211X1 U128 ( .C(n185), .D(n20), .A(n32), .B(n171), .Y(n144) );
  AND2X1 U129 ( .A(n140), .B(n132), .Y(n100) );
  OAI21X1 U130 ( .B(n22), .C(n189), .A(n177), .Y(n169) );
  NOR2X1 U131 ( .A(n137), .B(n138), .Y(n95) );
  OAI21X1 U132 ( .B(n176), .C(n23), .A(n180), .Y(n173) );
  NOR3XL U133 ( .A(n131), .B(n140), .C(n150), .Y(n182) );
  NAND2X1 U134 ( .A(n148), .B(n149), .Y(n113) );
  NAND2X1 U135 ( .A(n155), .B(n191), .Y(n187) );
  NAND2X1 U136 ( .A(n145), .B(n193), .Y(n161) );
  NOR2X1 U137 ( .A(n141), .B(n134), .Y(n103) );
  NAND2X1 U138 ( .A(n146), .B(n147), .Y(n94) );
  NOR32XL U139 ( .B(n179), .C(n137), .A(n162), .Y(n176) );
  NAND21X1 U140 ( .B(n138), .A(n162), .Y(n93) );
  NAND32X1 U141 ( .B(n163), .C(n146), .A(n172), .Y(n166) );
  AND2X1 U142 ( .A(n135), .B(n136), .Y(n127) );
  NOR3XL U143 ( .A(n165), .B(n148), .C(n164), .Y(n185) );
  NAND2X1 U144 ( .A(n150), .B(n132), .Y(n129) );
  NOR2X1 U145 ( .A(n156), .B(n134), .Y(n124) );
  NOR2X1 U146 ( .A(n185), .B(n27), .Y(n188) );
  NAND2X1 U147 ( .A(n163), .B(n147), .Y(n91) );
  NAND2X1 U148 ( .A(n164), .B(n149), .Y(n126) );
  NOR2X1 U149 ( .A(n133), .B(n134), .Y(n116) );
  NAND2X1 U150 ( .A(n131), .B(n132), .Y(n118) );
  NOR2X1 U151 ( .A(n135), .B(n139), .Y(n184) );
  ENOX1 U152 ( .A(n35), .B(n75), .C(n76), .D(intcall), .Y(int_ack_03) );
  OAI21X1 U153 ( .B(n39), .C(n37), .A(n60), .Y(n76) );
  AND3X1 U154 ( .A(n60), .B(n61), .C(n34), .Y(n55) );
  NOR2X1 U155 ( .A(n73), .B(n35), .Y(int_ack_43) );
  AOI211X1 U156 ( .C(n66), .D(n67), .A(int_ack_03), .B(int_ack_43), .Y(n50) );
  OAI32X1 U157 ( .A(n202), .B(n21), .C(n40), .D(n41), .E(n201), .Y(n196) );
  OA21X1 U158 ( .B(n42), .C(n43), .A(n44), .Y(n41) );
  OAI21X1 U159 ( .B(n45), .C(n44), .A(n46), .Y(n197) );
  GEN2XL U160 ( .D(n47), .E(n38), .C(n43), .B(n44), .A(n36), .Y(n46) );
  OAI31XL U161 ( .A(n45), .B(n40), .C(n202), .D(n49), .Y(n199) );
  GEN2XL U162 ( .D(n42), .E(n201), .C(n43), .B(n202), .A(n32), .Y(n49) );
  NAND2X1 U163 ( .A(n48), .B(n40), .Y(n44) );
  NOR21XL U164 ( .B(n62), .A(n63), .Y(n53) );
  NOR21XL U165 ( .B(n62), .A(n65), .Y(n56) );
  NOR21XL U166 ( .B(n62), .A(n64), .Y(n57) );
  NOR2X1 U167 ( .A(n65), .B(n75), .Y(int_ack_13) );
  AND2X1 U168 ( .A(n60), .B(n37), .Y(n62) );
  NOR2X1 U169 ( .A(n64), .B(n75), .Y(int_ack_0b) );
  NOR2X1 U170 ( .A(n63), .B(n73), .Y(int_ack_5b) );
  NOR2X1 U171 ( .A(n65), .B(n73), .Y(int_ack_53) );
  NOR2X1 U172 ( .A(n64), .B(n73), .Y(int_ack_4b) );
  NOR2X1 U173 ( .A(n34), .B(n72), .Y(int_ack_6b) );
  NOR2X1 U174 ( .A(n63), .B(n75), .Y(int_ack_1b) );
  OAI22X1 U175 ( .A(n47), .B(n38), .C(n21), .D(n44), .Y(n198) );
  INVX1 U176 ( .A(n45), .Y(n21) );
  INVX1 U177 ( .A(n66), .Y(n35) );
  NOR2X1 U178 ( .A(n65), .B(n33), .Y(int_ack_93) );
  NOR2X1 U179 ( .A(n64), .B(n33), .Y(int_ack_8b) );
  INVX1 U180 ( .A(n67), .Y(n33) );
  NOR21XL U181 ( .B(n147), .A(n172), .Y(n120) );
  AND2X1 U182 ( .A(n149), .B(n165), .Y(n122) );
  NOR2X1 U183 ( .A(n179), .B(n138), .Y(n115) );
  NOR3XL U184 ( .A(n71), .B(n37), .C(n35), .Y(int_ack_a3) );
  NOR3XL U185 ( .A(n71), .B(n37), .C(n64), .Y(int_ack_ab) );
  NOR2X1 U186 ( .A(n63), .B(n33), .Y(int_ack_9b) );
  AND2X1 U187 ( .A(irq_r), .B(ien0[7]), .Y(irq) );
  NOR21XL U188 ( .B(ien1[0]), .A(n195), .Y(n135) );
  AOI22X1 U189 ( .A(int_vect_43), .B(n31), .C(sdaiff), .D(isr_tm), .Y(n195) );
  NOR32XL U190 ( .B(ien1[2]), .C(int_vect_53), .A(n131), .Y(n150) );
  AOI21X1 U191 ( .B(n166), .C(ip0[4]), .A(n173), .Y(n171) );
  NAND32X1 U192 ( .B(n188), .C(is_reg[1]), .A(n170), .Y(n142) );
  NAND21X1 U193 ( .B(n182), .A(ip1[2]), .Y(n191) );
  OAI221X1 U194 ( .A(n24), .B(n151), .C(n152), .D(n29), .E(n153), .Y(n132) );
  INVX1 U195 ( .A(ip1[2]), .Y(n29) );
  AOI21X1 U196 ( .B(n154), .C(ip0[2]), .A(n155), .Y(n152) );
  OAI221X1 U197 ( .A(n22), .B(n173), .C(n174), .D(n28), .E(n167), .Y(n147) );
  INVX1 U198 ( .A(ip1[4]), .Y(n28) );
  AOI21X1 U199 ( .B(n177), .C(ip0[4]), .A(n178), .Y(n174) );
  AOI221XL U200 ( .A(ip0[1]), .B(n157), .C(n158), .D(ip1[1]), .E(n159), .Y(
        n134) );
  OAI21X1 U201 ( .B(n160), .C(n25), .A(n161), .Y(n158) );
  AND2X1 U202 ( .A(int_vect_93), .B(ien2[2]), .Y(n131) );
  NAND21X1 U203 ( .B(n183), .A(ip1[1]), .Y(n192) );
  AOI221XL U204 ( .A(ip0[3]), .B(n180), .C(n181), .D(ip1[3]), .E(n175), .Y(
        n138) );
  OAI21X1 U205 ( .B(n186), .C(n23), .A(n187), .Y(n181) );
  OAI211X1 U206 ( .C(n26), .D(n193), .A(n38), .B(ien0[7]), .Y(n160) );
  AND2X1 U207 ( .A(int_vect_03), .B(ien0[0]), .Y(n139) );
  OAI21X1 U208 ( .B(n139), .C(n135), .A(ip1[0]), .Y(n193) );
  AOI211X1 U209 ( .C(ip0[5]), .D(n188), .A(is_reg[2]), .B(n169), .Y(n145) );
  INVX1 U210 ( .A(isr_tm), .Y(n31) );
  NAND2X1 U211 ( .A(int_vect_8b), .B(ien2[1]), .Y(n133) );
  NAND4X1 U212 ( .A(int_vect_4b), .B(ien1[1]), .C(n133), .D(n31), .Y(n156) );
  NAND3X1 U213 ( .A(ien0[1]), .B(n31), .C(int_vect_0b), .Y(n141) );
  NOR21XL U214 ( .B(ien0[4]), .A(n194), .Y(n146) );
  AOI22X1 U215 ( .A(int_vect_23), .B(n31), .C(rxd0ff), .D(isr_tm), .Y(n194) );
  AND3X1 U216 ( .A(ien1[3]), .B(n179), .C(int_vect_5b), .Y(n162) );
  NAND21X1 U217 ( .B(n176), .A(ip1[3]), .Y(n190) );
  AND2X1 U218 ( .A(ien0[5]), .B(i2c_int), .Y(n148) );
  AND2X1 U219 ( .A(int_vect_13), .B(ien0[2]), .Y(n140) );
  OAI221X1 U220 ( .A(n26), .B(n142), .C(n143), .D(n30), .E(n144), .Y(n136) );
  AOI31X1 U221 ( .A(ip0[0]), .B(n38), .C(ien0[7]), .D(n145), .Y(n143) );
  INVX1 U222 ( .A(ip0[0]), .Y(n26) );
  INVX1 U223 ( .A(is_reg[3]), .Y(n38) );
  NAND3X1 U224 ( .A(ien0[3]), .B(n31), .C(int_vect_1b), .Y(n137) );
  NAND2X1 U225 ( .A(ip1[4]), .B(n166), .Y(n189) );
  NOR32XL U226 ( .B(ien1[5]), .C(int_vect_6b), .A(n165), .Y(n164) );
  AND3X1 U227 ( .A(ien1[4]), .B(n172), .C(int_vect_63), .Y(n163) );
  INVX1 U228 ( .A(ip0[2]), .Y(n24) );
  INVX1 U229 ( .A(ip0[3]), .Y(n23) );
  INVX1 U230 ( .A(ip0[1]), .Y(n25) );
  INVX1 U231 ( .A(ip1[5]), .Y(n27) );
  INVX1 U232 ( .A(ip0[4]), .Y(n22) );
  INVX1 U233 ( .A(ip0[5]), .Y(n20) );
  INVX1 U234 ( .A(is_reg[0]), .Y(n32) );
  INVX1 U235 ( .A(ip1[0]), .Y(n30) );
  NOR32XL U236 ( .B(n36), .C(n47), .A(is_reg[3]), .Y(n42) );
  NAND21X1 U237 ( .B(intvect[3]), .A(n74), .Y(n75) );
  OAI211X1 U238 ( .C(n50), .D(n30), .A(n51), .B(n52), .Y(n40) );
  AOI22X1 U239 ( .A(ip1[2]), .B(n56), .C(ip1[1]), .D(n57), .Y(n51) );
  AOI222XL U240 ( .A(ip1[3]), .B(n53), .C(ip1[5]), .D(n54), .E(ip1[4]), .F(n55), .Y(n52) );
  AND3X1 U241 ( .A(n61), .B(n60), .C(intvect[0]), .Y(n54) );
  NOR3XL U242 ( .A(intvect[2]), .B(intvect[4]), .C(n203), .Y(n74) );
  NOR3XL U243 ( .A(n203), .B(intvect[1]), .C(n37), .Y(n61) );
  NAND2X1 U244 ( .A(n74), .B(intvect[3]), .Y(n73) );
  NAND31X1 U245 ( .C(intvect[4]), .A(intvect[3]), .B(n61), .Y(n72) );
  NAND31X1 U246 ( .C(intvect[3]), .A(intcall), .B(intvect[4]), .Y(n71) );
  OAI211X1 U247 ( .C(n50), .D(n26), .A(n58), .B(n59), .Y(n45) );
  AOI22X1 U248 ( .A(ip0[2]), .B(n56), .C(ip0[1]), .D(n57), .Y(n58) );
  AOI222XL U249 ( .A(ip0[3]), .B(n53), .C(ip0[5]), .D(n54), .E(ip0[4]), .F(n55), .Y(n59) );
  NOR2X1 U250 ( .A(intvect[0]), .B(n72), .Y(int_ack_63) );
  NOR2X1 U251 ( .A(n71), .B(intvect[2]), .Y(n67) );
  NOR2X1 U252 ( .A(intvect[0]), .B(intvect[1]), .Y(n66) );
  INVX1 U253 ( .A(intvect[0]), .Y(n34) );
  INVX1 U254 ( .A(intvect[1]), .Y(n39) );
  INVX1 U255 ( .A(intvect[2]), .Y(n37) );
  NAND2X1 U256 ( .A(intvect[4]), .B(intvect[3]), .Y(n60) );
  NAND2X1 U257 ( .A(intvect[0]), .B(n39), .Y(n64) );
  NAND2X1 U258 ( .A(intvect[1]), .B(intvect[0]), .Y(n63) );
  NAND2X1 U259 ( .A(intvect[1]), .B(n34), .Y(n65) );
  INVX1 U260 ( .A(is_reg[2]), .Y(n36) );
  INVX1 U261 ( .A(is_reg[1]), .Y(n201) );
  AND2X1 U262 ( .A(int_vect_ab), .B(ien2[5]), .Y(n165) );
  NAND2X1 U263 ( .A(int_vect_a3), .B(ien2[4]), .Y(n172) );
  NAND2X1 U264 ( .A(int_vect_9b), .B(ien2[3]), .Y(n179) );
endmodule


module SNPS_CLOCK_GATE_HIGH_isr_a0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_isr_a0_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_isr_a0_3 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_isr_a0_4 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_isr_a0_5 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_isr_a0_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module watchdog_a0 ( wdt_slow, clkwdt, clkper, resetff, newinstr, wdts_s, wdts, 
        ip0wdts, wdt_tm, sfrdatai, sfraddr, sfrwe, wdtrel );
  output [1:0] wdts_s;
  input [7:0] sfrdatai;
  input [6:0] sfraddr;
  output [7:0] wdtrel;
  input wdt_slow, clkwdt, clkper, resetff, newinstr, sfrwe;
  output wdts, ip0wdts, wdt_tm;
  wire   wdt_tm_sync, wdt_act_sync, wdt_act, wdtrefresh_sync, N26, N27, N28,
         N29, N30, N31, N32, N33, N34, N67, N68, N69, N70, N71, pres_2, N112,
         N113, N114, N115, N116, N130, N131, N132, N133, N134, N135, N136,
         N137, N138, N139, N140, N141, N142, N143, N144, N165, N166, N167,
         N168, N169, N170, N171, N172, N173, N174, N175, N176, N177, N178,
         N179, N180, wdt_normal, wdt_normal_ff, N212, net12155, net12161,
         net12166, net12171, net12176, n21, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, add_93_carry_2_,
         add_93_carry_3_, add_93_carry_4_, add_93_carry_5_, add_93_carry_6_,
         n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n22, n23, n24;
  wire   [14:9] half_RSL_tmp;
  wire   [1:0] pres_8;
  wire   [3:0] cycles_reg;
  wire   [3:0] pres_16;
  wire   [6:0] wdth;
  wire   [7:0] wdtl;

  SNPS_CLOCK_GATE_HIGH_watchdog_a0_0 clk_gate_wdtrel_s_reg ( .CLK(clkper), 
        .EN(N26), .ENCLK(net12155), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_watchdog_a0_4 clk_gate_cycles_reg_reg ( .CLK(clkwdt), 
        .EN(N67), .ENCLK(net12161), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_watchdog_a0_3 clk_gate_pres_16_reg ( .CLK(clkwdt), .EN(
        N112), .ENCLK(net12166), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_watchdog_a0_2 clk_gate_wdth_reg ( .CLK(clkwdt), .EN(
        N165), .ENCLK(net12171), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_watchdog_a0_1 clk_gate_wdtl_reg ( .CLK(clkwdt), .EN(n21), .ENCLK(net12176), .TE(1'b0) );
  watchdog_a0_DW01_inc_0 add_278 ( .A(wdtl), .SUM({N144, N143, N142, N141, 
        N140, N139, N138, N137}) );
  watchdog_a0_DW01_inc_1 add_272 ( .A(wdth), .SUM({N136, N135, N134, N133, 
        N132, N131, N130}) );
  DFFQX1 wdts_s_reg_1_ ( .D(n126), .C(net12176), .Q(wdts_s[1]) );
  DFFQX1 wdt_act_reg ( .D(n130), .C(clkper), .Q(wdt_act) );
  DFFQX1 wdts_reg ( .D(wdts_s[0]), .C(clkper), .Q(wdts) );
  DFFQX1 wdt_normal_ff_reg ( .D(n3), .C(clkper), .Q(wdt_normal_ff) );
  DFFQX1 pres_2_reg ( .D(n127), .C(net12161), .Q(pres_2) );
  DFFQX1 wdt_tm_sync_reg ( .D(wdt_tm), .C(clkwdt), .Q(wdt_tm_sync) );
  DFFQX1 wdt_normal_reg ( .D(n133), .C(clkper), .Q(wdt_normal) );
  DFFQX1 wdts_s_reg_0_ ( .D(n132), .C(net12176), .Q(wdts_s[0]) );
  DFFQX1 wdt_act_sync_reg ( .D(wdt_act), .C(clkwdt), .Q(wdt_act_sync) );
  DFFQX1 pres_16_reg_3_ ( .D(N116), .C(net12166), .Q(pres_16[3]) );
  DFFQX1 wdth_reg_6_ ( .D(N172), .C(net12171), .Q(wdth[6]) );
  DFFQX1 pres_8_reg_0_ ( .D(n129), .C(net12161), .Q(pres_8[0]) );
  DFFQX1 pres_8_reg_1_ ( .D(n128), .C(net12161), .Q(pres_8[1]) );
  DFFQX1 wdtl_reg_2_ ( .D(N175), .C(net12176), .Q(wdtl[2]) );
  DFFQX1 wdtrefresh_reg ( .D(N212), .C(clkper), .Q(wdtrefresh_sync) );
  DFFQX1 cycles_reg_reg_2_ ( .D(N70), .C(net12161), .Q(cycles_reg[2]) );
  DFFQX1 pres_16_reg_1_ ( .D(N114), .C(net12166), .Q(pres_16[1]) );
  DFFQX1 cycles_reg_reg_1_ ( .D(N69), .C(net12161), .Q(cycles_reg[1]) );
  DFFQX1 wdtl_reg_1_ ( .D(N174), .C(net12176), .Q(wdtl[1]) );
  DFFQX1 wdtl_reg_7_ ( .D(N180), .C(net12176), .Q(wdtl[7]) );
  DFFQX1 wdtl_reg_0_ ( .D(N173), .C(net12176), .Q(wdtl[0]) );
  DFFQX1 pres_16_reg_0_ ( .D(N113), .C(net12166), .Q(pres_16[0]) );
  DFFQX1 cycles_reg_reg_0_ ( .D(N68), .C(net12161), .Q(cycles_reg[0]) );
  DFFQX1 wdth_reg_1_ ( .D(N167), .C(net12171), .Q(wdth[1]) );
  DFFQX1 wdth_reg_3_ ( .D(N169), .C(net12171), .Q(wdth[3]) );
  DFFQX1 wdth_reg_0_ ( .D(N166), .C(net12171), .Q(wdth[0]) );
  DFFQX1 wdtl_reg_3_ ( .D(N176), .C(net12176), .Q(wdtl[3]) );
  DFFQX1 wdth_reg_2_ ( .D(N168), .C(net12171), .Q(wdth[2]) );
  DFFQX1 pres_16_reg_2_ ( .D(N115), .C(net12166), .Q(pres_16[2]) );
  DFFQX1 cycles_reg_reg_3_ ( .D(N71), .C(net12161), .Q(cycles_reg[3]) );
  DFFQX1 wdtl_reg_4_ ( .D(N177), .C(net12176), .Q(wdtl[4]) );
  DFFQX1 wdth_reg_4_ ( .D(N170), .C(net12171), .Q(wdth[4]) );
  DFFQX1 wdth_reg_5_ ( .D(N171), .C(net12171), .Q(wdth[5]) );
  DFFQX1 wdtl_reg_5_ ( .D(N178), .C(net12176), .Q(wdtl[5]) );
  DFFQX1 wdtl_reg_6_ ( .D(N179), .C(net12176), .Q(wdtl[6]) );
  DFFQX1 wdtrel_s_reg_7_ ( .D(N34), .C(net12155), .Q(wdtrel[7]) );
  DFFQX1 ip0wdts_reg ( .D(n131), .C(clkper), .Q(ip0wdts) );
  DFFQX1 wdtrel_s_reg_6_ ( .D(N33), .C(net12155), .Q(wdtrel[6]) );
  DFFQX1 wdtrel_s_reg_3_ ( .D(N30), .C(net12155), .Q(wdtrel[3]) );
  DFFQX1 wdtrel_s_reg_1_ ( .D(N28), .C(net12155), .Q(wdtrel[1]) );
  DFFQX1 wdtrel_s_reg_2_ ( .D(N29), .C(net12155), .Q(wdtrel[2]) );
  DFFQX1 wdt_tm_s_reg ( .D(n134), .C(clkper), .Q(wdt_tm) );
  DFFQX1 wdtrel_s_reg_5_ ( .D(N32), .C(net12155), .Q(wdtrel[5]) );
  DFFQX1 wdtrel_s_reg_4_ ( .D(N31), .C(net12155), .Q(wdtrel[4]) );
  DFFQX1 wdtrel_s_reg_0_ ( .D(N27), .C(net12155), .Q(wdtrel[0]) );
  BUFX2 U3 ( .A(resetff), .Y(n1) );
  NAND32XL U4 ( .B(sfraddr[4]), .C(sfraddr[6]), .A(sfrwe), .Y(n95) );
  NAND4XL U5 ( .A(sfraddr[1]), .B(n5), .C(sfraddr[2]), .D(n106), .Y(n105) );
  INVX1 U6 ( .A(n95), .Y(n5) );
  NOR43XL U7 ( .B(n107), .C(n108), .D(sfraddr[3]), .A(sfraddr[0]), .Y(n77) );
  NOR3XL U8 ( .A(sfraddr[1]), .B(sfraddr[6]), .C(sfraddr[2]), .Y(n107) );
  AND4X1 U9 ( .A(sfraddr[4]), .B(sfraddr[5]), .C(sfrwe), .D(sfrdatai[6]), .Y(
        n108) );
  INVX1 U10 ( .A(n89), .Y(n4) );
  NAND4X1 U11 ( .A(sfraddr[5]), .B(sfraddr[3]), .C(n5), .D(n91), .Y(n90) );
  NOR3XL U12 ( .A(sfraddr[0]), .B(sfraddr[2]), .C(sfraddr[1]), .Y(n91) );
  NOR31X1 U13 ( .C(sfraddr[3]), .A(sfraddr[2]), .B(sfraddr[1]), .Y(n81) );
  INVX1 U14 ( .A(sfrdatai[6]), .Y(n2) );
  NAND2X1 U15 ( .A(n69), .B(n12), .Y(n121) );
  NOR32XL U16 ( .B(n23), .C(n90), .A(newinstr), .Y(n89) );
  NOR21XL U17 ( .B(sfrdatai[0]), .A(n105), .Y(N27) );
  NOR21XL U18 ( .B(sfrdatai[1]), .A(n105), .Y(N28) );
  NOR21XL U19 ( .B(sfrdatai[2]), .A(n105), .Y(N29) );
  NOR21XL U20 ( .B(sfrdatai[3]), .A(n105), .Y(N30) );
  NOR21XL U21 ( .B(sfrdatai[4]), .A(n105), .Y(N31) );
  NOR21XL U22 ( .B(sfrdatai[5]), .A(n105), .Y(N32) );
  NOR21XL U23 ( .B(sfrdatai[7]), .A(n105), .Y(N34) );
  NOR2X1 U24 ( .A(n2), .B(n105), .Y(N33) );
  NAND2X1 U25 ( .A(n23), .B(n105), .Y(N26) );
  NOR3XL U26 ( .A(n49), .B(n22), .C(n20), .Y(n85) );
  NAND2X1 U27 ( .A(n110), .B(n50), .Y(n43) );
  AND2X1 U28 ( .A(n73), .B(n115), .Y(n69) );
  OAI21X1 U29 ( .B(n123), .C(n121), .A(n103), .Y(N115) );
  XNOR2XL U30 ( .A(n122), .B(n10), .Y(n123) );
  NOR2X1 U31 ( .A(n10), .B(n122), .Y(n116) );
  OAI211X1 U32 ( .C(n50), .D(n113), .A(n8), .B(n23), .Y(N165) );
  INVX1 U33 ( .A(n112), .Y(n8) );
  NAND2X1 U34 ( .A(n111), .B(n110), .Y(n113) );
  NOR21XL U35 ( .B(N143), .A(n43), .Y(N179) );
  NOR21XL U36 ( .B(N142), .A(n43), .Y(N178) );
  NOR21XL U37 ( .B(N141), .A(n43), .Y(N177) );
  NOR21XL U38 ( .B(N140), .A(n43), .Y(N176) );
  NOR21XL U39 ( .B(N139), .A(n43), .Y(N175) );
  NOR21XL U40 ( .B(N138), .A(n43), .Y(N174) );
  INVX1 U41 ( .A(n72), .Y(n12) );
  NOR2X1 U42 ( .A(n16), .B(n15), .Y(n115) );
  NAND2X1 U43 ( .A(n99), .B(n12), .Y(n96) );
  INVX1 U44 ( .A(n101), .Y(n13) );
  NAND2X1 U45 ( .A(n23), .B(n72), .Y(N67) );
  OAI32X1 U46 ( .A(n90), .B(resetff), .C(n2), .D(n7), .E(n4), .Y(n133) );
  INVX1 U47 ( .A(wdt_normal), .Y(n7) );
  OAI21X1 U48 ( .B(n2), .C(n92), .A(n93), .Y(n134) );
  NAND3X1 U49 ( .A(n92), .B(n23), .C(wdt_tm), .Y(n93) );
  NAND4XL U50 ( .A(sfraddr[1]), .B(sfraddr[0]), .C(sfraddr[2]), .D(n94), .Y(
        n92) );
  NOR4XL U51 ( .A(sfraddr[5]), .B(sfraddr[3]), .C(resetff), .D(n95), .Y(n94)
         );
  ENOX1 U52 ( .A(n1), .B(n76), .C(wdt_act), .D(n76), .Y(n130) );
  OAI21X1 U53 ( .B(n77), .C(resetff), .A(n11), .Y(n76) );
  INVX1 U54 ( .A(n88), .Y(n3) );
  AOI32X1 U55 ( .A(wdt_normal), .B(n23), .C(n4), .D(n89), .E(wdt_normal_ff), 
        .Y(n88) );
  NOR4XL U56 ( .A(sfraddr[5]), .B(sfraddr[3]), .C(sfraddr[0]), .D(resetff), 
        .Y(n106) );
  AND3X1 U57 ( .A(n77), .B(wdt_normal_ff), .C(n23), .Y(N212) );
  OAI21X1 U58 ( .B(n1), .C(n78), .A(n79), .Y(n131) );
  NAND3X1 U59 ( .A(n80), .B(n23), .C(ip0wdts), .Y(n79) );
  EORX1 U60 ( .A(wdts_s[0]), .B(n80), .C(n80), .D(n2), .Y(n78) );
  NAND4X1 U61 ( .A(n5), .B(sfraddr[5]), .C(sfraddr[0]), .D(n81), .Y(n80) );
  XNOR2XL U62 ( .A(half_RSL_tmp[14]), .B(n22), .Y(n56) );
  OAI21X1 U63 ( .B(n43), .C(n44), .A(n45), .Y(n126) );
  NAND41X1 U64 ( .D(n46), .A(wdts_s[1]), .B(n47), .C(n44), .Y(n45) );
  OAI31XL U65 ( .A(n18), .B(n48), .C(n49), .D(n50), .Y(n46) );
  NAND3X1 U66 ( .A(n51), .B(n52), .C(n53), .Y(n44) );
  NOR4XL U67 ( .A(n54), .B(n55), .C(n56), .D(n57), .Y(n53) );
  XOR2X1 U68 ( .A(n58), .B(wdtl[7]), .Y(n55) );
  NAND4X1 U69 ( .A(n59), .B(n60), .C(n61), .D(n62), .Y(n54) );
  XNOR2XL U70 ( .A(half_RSL_tmp[13]), .B(n20), .Y(n57) );
  XNOR2XL U71 ( .A(wdth[2]), .B(half_RSL_tmp[11]), .Y(n62) );
  XNOR2XL U72 ( .A(wdth[3]), .B(half_RSL_tmp[12]), .Y(n59) );
  XNOR2XL U73 ( .A(wdth[1]), .B(half_RSL_tmp[10]), .Y(n61) );
  XNOR2XL U74 ( .A(wdth[0]), .B(half_RSL_tmp[9]), .Y(n60) );
  OAI22AX1 U75 ( .D(n82), .C(n43), .A(n11), .B(n82), .Y(n132) );
  OAI211X1 U76 ( .C(n83), .D(n84), .A(n50), .B(n47), .Y(n82) );
  NAND4X1 U77 ( .A(n86), .B(n18), .C(wdth[2]), .D(n87), .Y(n83) );
  NAND3X1 U78 ( .A(n48), .B(wdth[6]), .C(n85), .Y(n84) );
  NAND4X1 U79 ( .A(n117), .B(n118), .C(wdtl[3]), .D(n119), .Y(n49) );
  AND2X1 U80 ( .A(wdtl[0]), .B(wdtl[1]), .Y(n119) );
  XNOR2XL U81 ( .A(n24), .B(wdtl[5]), .Y(n117) );
  XNOR2XL U82 ( .A(n24), .B(wdtl[6]), .Y(n118) );
  NAND42X1 U83 ( .C(n49), .D(n18), .A(wdtl[4]), .B(n86), .Y(n50) );
  NOR43XL U84 ( .B(n114), .C(n115), .D(n104), .A(n17), .Y(n111) );
  OAI21BBX1 U85 ( .A(n116), .B(pres_16[3]), .C(wdtrel[7]), .Y(n114) );
  NOR21XL U86 ( .B(n104), .A(wdtrefresh_sync), .Y(n73) );
  NOR21XL U87 ( .B(N144), .A(n43), .Y(N180) );
  XNOR2XL U88 ( .A(wdtl[4]), .B(wdt_slow), .Y(n48) );
  NAND32X1 U89 ( .B(n73), .C(wdt_tm_sync), .A(n47), .Y(n70) );
  AO22X1 U90 ( .A(wdtrel[6]), .B(n112), .C(N136), .D(n110), .Y(N172) );
  NAND2X1 U91 ( .A(cycles_reg[1]), .B(cycles_reg[0]), .Y(n101) );
  NOR3XL U92 ( .A(n101), .B(cycles_reg[2]), .C(n14), .Y(n104) );
  NOR42XL U93 ( .C(wdtl[2]), .D(wdtl[0]), .A(n64), .B(n65), .Y(n51) );
  XOR2X1 U94 ( .A(n66), .B(wdtl[4]), .Y(n64) );
  XNOR2XL U95 ( .A(n24), .B(wdtl[3]), .Y(n65) );
  NAND2X1 U96 ( .A(wdt_slow), .B(wdtrel[0]), .Y(n66) );
  OAI31XL U97 ( .A(n96), .B(n13), .C(n14), .D(n97), .Y(N71) );
  OAI21X1 U98 ( .B(n98), .C(wdt_tm_sync), .A(n12), .Y(n97) );
  AND4X1 U99 ( .A(n14), .B(cycles_reg[2]), .C(n99), .D(n13), .Y(n98) );
  AOI211X1 U100 ( .C(n24), .D(n19), .A(n63), .B(wdtl[1]), .Y(n52) );
  ENOX1 U101 ( .A(wdtl[5]), .B(n19), .C(wdt_slow), .D(wdtl[5]), .Y(n63) );
  INVX1 U102 ( .A(wdtl[6]), .Y(n19) );
  OAI21X1 U103 ( .B(n120), .C(n121), .A(n103), .Y(N116) );
  XNOR2XL U104 ( .A(pres_16[3]), .B(n116), .Y(n120) );
  OAI21X1 U105 ( .B(n124), .C(n121), .A(n103), .Y(N114) );
  XNOR2XL U106 ( .A(pres_16[1]), .B(pres_16[0]), .Y(n124) );
  OAI21X1 U107 ( .B(pres_16[0]), .C(n121), .A(n103), .Y(N113) );
  NOR2X1 U108 ( .A(n104), .B(wdtrefresh_sync), .Y(n99) );
  OAI22X1 U109 ( .A(n15), .B(n70), .C(n75), .D(n72), .Y(n129) );
  AOI21X1 U110 ( .B(n73), .C(n15), .A(wdt_tm_sync), .Y(n75) );
  OAI22X1 U111 ( .A(n16), .B(n70), .C(n71), .D(n72), .Y(n128) );
  AOI21X1 U112 ( .B(n73), .C(n74), .A(wdt_tm_sync), .Y(n71) );
  XNOR2XL U113 ( .A(n15), .B(pres_8[1]), .Y(n74) );
  OAI32X1 U114 ( .A(n67), .B(resetff), .C(n6), .D(n68), .E(n17), .Y(n127) );
  AOI21X1 U115 ( .B(n17), .C(n9), .A(wdt_tm_sync), .Y(n67) );
  INVX1 U116 ( .A(n68), .Y(n6) );
  NAND32X1 U117 ( .B(n69), .C(wdt_tm_sync), .A(n47), .Y(n68) );
  NAND2X1 U118 ( .A(pres_16[1]), .B(pres_16[0]), .Y(n122) );
  OAI211X1 U119 ( .C(n125), .D(n72), .A(n103), .B(n23), .Y(N112) );
  AOI21X1 U120 ( .B(n69), .C(pres_2), .A(wdtrefresh_sync), .Y(n125) );
  NOR2X1 U121 ( .A(wdt_slow), .B(wdtrel[0]), .Y(n58) );
  INVX1 U122 ( .A(wdth[4]), .Y(n20) );
  INVX1 U123 ( .A(wdth[5]), .Y(n22) );
  INVX1 U124 ( .A(pres_16[2]), .Y(n10) );
  INVX1 U125 ( .A(cycles_reg[3]), .Y(n14) );
  INVX1 U126 ( .A(n109), .Y(n21) );
  AOI211X1 U127 ( .C(n110), .D(n111), .A(n112), .B(resetff), .Y(n109) );
  XNOR2XL U128 ( .A(wdtl[7]), .B(n24), .Y(n86) );
  NOR21XL U129 ( .B(N137), .A(n43), .Y(N173) );
  INVX1 U130 ( .A(resetff), .Y(n23) );
  NOR2X1 U131 ( .A(n9), .B(resetff), .Y(n112) );
  NAND2X1 U132 ( .A(wdt_act_sync), .B(n23), .Y(n72) );
  AO22X1 U133 ( .A(wdtrel[5]), .B(n112), .C(N135), .D(n110), .Y(N171) );
  AO22X1 U134 ( .A(wdtrel[4]), .B(n112), .C(N134), .D(n110), .Y(N170) );
  AO22X1 U135 ( .A(wdtrel[3]), .B(n112), .C(N133), .D(n110), .Y(N169) );
  AO22X1 U136 ( .A(wdtrel[2]), .B(n112), .C(N132), .D(n110), .Y(N168) );
  AO22X1 U137 ( .A(wdtrel[1]), .B(n112), .C(N131), .D(n110), .Y(N167) );
  AO22X1 U138 ( .A(wdtrel[0]), .B(n112), .C(N130), .D(n110), .Y(N166) );
  NOR2X1 U139 ( .A(n72), .B(wdtrefresh_sync), .Y(n110) );
  AND3X1 U140 ( .A(wdth[3]), .B(wdth[1]), .C(wdth[0]), .Y(n87) );
  NOR2X1 U141 ( .A(wdtrefresh_sync), .B(resetff), .Y(n47) );
  NAND2X1 U142 ( .A(wdt_tm_sync), .B(n12), .Y(n103) );
  OAI21X1 U143 ( .B(n102), .C(n96), .A(n103), .Y(N69) );
  XNOR2XL U144 ( .A(cycles_reg[1]), .B(cycles_reg[0]), .Y(n102) );
  OAI21X1 U145 ( .B(cycles_reg[0]), .C(n96), .A(n103), .Y(N68) );
  INVX1 U146 ( .A(pres_8[0]), .Y(n15) );
  INVX1 U147 ( .A(wdtl[2]), .Y(n18) );
  NOR3XL U148 ( .A(n96), .B(wdt_tm_sync), .C(n100), .Y(N70) );
  XNOR2XL U149 ( .A(n13), .B(cycles_reg[2]), .Y(n100) );
  INVX1 U150 ( .A(pres_8[1]), .Y(n16) );
  INVX1 U151 ( .A(wdtrefresh_sync), .Y(n9) );
  INVX1 U152 ( .A(pres_2), .Y(n17) );
  INVX1 U153 ( .A(wdts_s[0]), .Y(n11) );
  INVX1 U154 ( .A(wdt_slow), .Y(n24) );
  XNOR2XL U155 ( .A(wdtrel[6]), .B(add_93_carry_6_), .Y(half_RSL_tmp[14]) );
  OR2X1 U156 ( .A(add_93_carry_5_), .B(wdtrel[5]), .Y(add_93_carry_6_) );
  XNOR2XL U157 ( .A(add_93_carry_5_), .B(wdtrel[5]), .Y(half_RSL_tmp[13]) );
  OR2X1 U158 ( .A(add_93_carry_4_), .B(wdtrel[4]), .Y(add_93_carry_5_) );
  XNOR2XL U159 ( .A(add_93_carry_4_), .B(wdtrel[4]), .Y(half_RSL_tmp[12]) );
  OR2X1 U160 ( .A(add_93_carry_3_), .B(wdtrel[3]), .Y(add_93_carry_4_) );
  XNOR2XL U161 ( .A(add_93_carry_3_), .B(wdtrel[3]), .Y(half_RSL_tmp[11]) );
  OR2X1 U162 ( .A(add_93_carry_2_), .B(wdtrel[2]), .Y(add_93_carry_3_) );
  XNOR2XL U163 ( .A(add_93_carry_2_), .B(wdtrel[2]), .Y(half_RSL_tmp[10]) );
  OR2X1 U164 ( .A(wdtrel[0]), .B(wdtrel[1]), .Y(add_93_carry_2_) );
  XNOR2XL U165 ( .A(wdtrel[0]), .B(wdtrel[1]), .Y(half_RSL_tmp[9]) );
endmodule


module watchdog_a0_DW01_inc_1 ( A, SUM );
  input [6:0] A;
  output [6:0] SUM;

  wire   [6:2] carry;

  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  XOR2X1 U1 ( .A(carry[6]), .B(A[6]), .Y(SUM[6]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module watchdog_a0_DW01_inc_0 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  XOR2X1 U1 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_watchdog_a0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_watchdog_a0_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_watchdog_a0_3 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_watchdog_a0_4 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_watchdog_a0_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module timer1_a0 ( clkper, rst, newinstr, t1ff, t1ack, int1ff, t1_tf1, t1ov, 
        sfrdatai, sfraddr, sfrwe, t1_tmod, t1_tr1, tl1, th1 );
  input [7:0] sfrdatai;
  input [6:0] sfraddr;
  output [3:0] t1_tmod;
  output [7:0] tl1;
  output [7:0] th1;
  input clkper, rst, newinstr, t1ff, t1ack, int1ff, sfrwe;
  output t1_tf1, t1ov, t1_tr1;
  wire   t1clr, th1_ov_ff, tl1_ov_ff, N31, N32, N33, N34, N35, N36, N37, N42,
         N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56,
         N57, N58, N68, N69, N70, N71, N72, N73, N74, N75, N76, N77, N78, N79,
         N80, N81, N82, N83, N84, N95, N96, N97, N98, clk_ov12, N100, net12193,
         net12199, net12204, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n59;
  wire   [1:0] t0_mode;
  wire   [3:0] clk_count;

  SNPS_CLOCK_GATE_HIGH_timer1_a0_0 clk_gate_t1_mode_reg ( .CLK(clkper), .EN(
        N31), .ENCLK(net12193), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_timer1_a0_2 clk_gate_tl1_s_reg ( .CLK(clkper), .EN(N50), 
        .ENCLK(net12199), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_timer1_a0_1 clk_gate_th1_s_reg ( .CLK(clkper), .EN(N76), 
        .ENCLK(net12204), .TE(1'b0) );
  timer1_a0_DW01_inc_0 add_278 ( .A(th1), .SUM({N75, N74, N73, N72, N71, N70, 
        N69, N68}) );
  timer1_a0_DW01_inc_1 add_244 ( .A(tl1), .SUM({N49, N48, N47, N46, N45, N44, 
        N43, N42}) );
  DFFQX1 th1_ov_ff_reg ( .D(n55), .C(clkper), .Q(th1_ov_ff) );
  DFFQX1 clk_count_reg_1_ ( .D(N96), .C(clkper), .Q(clk_count[1]) );
  DFFQX1 clk_count_reg_2_ ( .D(N97), .C(clkper), .Q(clk_count[2]) );
  DFFQX1 clk_count_reg_0_ ( .D(N95), .C(clkper), .Q(clk_count[0]) );
  DFFQX1 clk_count_reg_3_ ( .D(N98), .C(clkper), .Q(clk_count[3]) );
  DFFQX1 t1clr_reg ( .D(n57), .C(clkper), .Q(t1clr) );
  DFFQX1 tl1_ov_ff_reg ( .D(n56), .C(clkper), .Q(tl1_ov_ff) );
  DFFQX1 clk_ov12_reg ( .D(N100), .C(clkper), .Q(clk_ov12) );
  DFFQX1 t0_mode_reg_1_ ( .D(N37), .C(net12193), .Q(t0_mode[1]) );
  DFFQX1 t0_mode_reg_0_ ( .D(N36), .C(net12193), .Q(t0_mode[0]) );
  DFFQX1 t1_ct_reg ( .D(N33), .C(net12193), .Q(t1_tmod[2]) );
  DFFQX1 t1_gate_reg ( .D(N32), .C(net12193), .Q(t1_tmod[3]) );
  DFFQX1 tl1_s_reg_7_ ( .D(N58), .C(net12199), .Q(tl1[7]) );
  DFFQX1 tl1_s_reg_5_ ( .D(N56), .C(net12199), .Q(tl1[5]) );
  DFFQX1 tl1_s_reg_6_ ( .D(N57), .C(net12199), .Q(tl1[6]) );
  DFFQX1 tl1_s_reg_1_ ( .D(N52), .C(net12199), .Q(tl1[1]) );
  DFFQX1 tl1_s_reg_3_ ( .D(N54), .C(net12199), .Q(tl1[3]) );
  DFFQX1 th1_s_reg_1_ ( .D(N78), .C(net12204), .Q(th1[1]) );
  DFFQX1 tl1_s_reg_2_ ( .D(N53), .C(net12199), .Q(tl1[2]) );
  DFFQX1 th1_s_reg_3_ ( .D(N80), .C(net12204), .Q(th1[3]) );
  DFFQX1 th1_s_reg_2_ ( .D(N79), .C(net12204), .Q(th1[2]) );
  DFFQX1 t1_tf1_s_reg ( .D(n54), .C(clkper), .Q(t1_tf1) );
  DFFQX1 th1_s_reg_7_ ( .D(N84), .C(net12204), .Q(th1[7]) );
  DFFQX1 tl1_s_reg_0_ ( .D(N51), .C(net12199), .Q(tl1[0]) );
  DFFQX1 th1_s_reg_5_ ( .D(N82), .C(net12204), .Q(th1[5]) );
  DFFQX1 th1_s_reg_4_ ( .D(N81), .C(net12204), .Q(th1[4]) );
  DFFQX1 tl1_s_reg_4_ ( .D(N55), .C(net12199), .Q(tl1[4]) );
  DFFQX1 th1_s_reg_0_ ( .D(N77), .C(net12204), .Q(th1[0]) );
  DFFQX1 t1_tr1_s_reg ( .D(n58), .C(clkper), .Q(t1_tr1) );
  DFFQX1 t1_mode_reg_0_ ( .D(N34), .C(net12193), .Q(t1_tmod[0]) );
  DFFQX1 t1_mode_reg_1_ ( .D(N35), .C(net12193), .Q(t1_tmod[1]) );
  DFFQX1 th1_s_reg_6_ ( .D(N83), .C(net12204), .Q(th1[6]) );
  NAND4XL U3 ( .A(sfraddr[2]), .B(sfraddr[0]), .C(n42), .D(n1), .Y(n41) );
  NAND21X1 U4 ( .B(n41), .A(n9), .Y(n39) );
  NAND2X1 U5 ( .A(n9), .B(n52), .Y(N31) );
  NOR21XL U6 ( .B(n42), .A(sfraddr[2]), .Y(n33) );
  NAND31X1 U7 ( .C(sfraddr[0]), .A(n1), .B(n33), .Y(n20) );
  NOR3XL U8 ( .A(n10), .B(rst), .C(n12), .Y(n43) );
  NOR2X1 U9 ( .A(n46), .B(n8), .Y(n45) );
  INVX1 U10 ( .A(n46), .Y(n10) );
  NAND4X1 U11 ( .A(sfraddr[0]), .B(n33), .C(n9), .D(n1), .Y(n52) );
  NOR2X1 U12 ( .A(n6), .B(n52), .Y(N33) );
  NOR2X1 U13 ( .A(n7), .B(n52), .Y(N32) );
  NOR2X1 U14 ( .A(n2), .B(n52), .Y(N36) );
  NOR2X1 U15 ( .A(n3), .B(n52), .Y(N37) );
  NOR2X1 U16 ( .A(n4), .B(n52), .Y(N34) );
  NOR2X1 U17 ( .A(n5), .B(n52), .Y(N35) );
  AND3X1 U18 ( .A(sfrwe), .B(sfraddr[3]), .C(n53), .Y(n42) );
  NOR3XL U19 ( .A(sfraddr[4]), .B(sfraddr[6]), .C(sfraddr[5]), .Y(n53) );
  OR4X1 U20 ( .A(n44), .B(n43), .C(n45), .D(n8), .Y(N50) );
  NAND3X1 U21 ( .A(sfraddr[0]), .B(n33), .C(sfraddr[1]), .Y(n46) );
  INVX1 U22 ( .A(n40), .Y(n11) );
  NAND3X1 U23 ( .A(n39), .B(n9), .C(n40), .Y(N76) );
  INVX1 U24 ( .A(sfraddr[1]), .Y(n1) );
  INVX1 U25 ( .A(sfrdatai[7]), .Y(n7) );
  INVX1 U26 ( .A(sfrdatai[0]), .Y(n2) );
  INVX1 U27 ( .A(sfrdatai[1]), .Y(n3) );
  INVX1 U28 ( .A(sfrdatai[4]), .Y(n4) );
  INVX1 U29 ( .A(sfrdatai[5]), .Y(n5) );
  INVX1 U30 ( .A(sfrdatai[6]), .Y(n6) );
  INVX1 U31 ( .A(n47), .Y(n12) );
  INVX1 U32 ( .A(n9), .Y(n8) );
  INVX1 U33 ( .A(rst), .Y(n9) );
  NOR4XL U34 ( .A(n48), .B(n47), .C(n10), .D(n8), .Y(n44) );
  AO22AXL U35 ( .A(N71), .B(n11), .C(sfrdatai[3]), .D(n39), .Y(N80) );
  AO22AXL U36 ( .A(N70), .B(n11), .C(sfrdatai[2]), .D(n39), .Y(N79) );
  NAND3X1 U37 ( .A(n41), .B(n9), .C(n30), .Y(n40) );
  ENOX1 U38 ( .A(n39), .B(n5), .C(N73), .D(n11), .Y(N82) );
  ENOX1 U39 ( .A(n39), .B(n4), .C(N72), .D(n11), .Y(N81) );
  ENOX1 U40 ( .A(n39), .B(n3), .C(N69), .D(n11), .Y(N78) );
  ENOX1 U41 ( .A(n6), .B(n39), .C(N74), .D(n11), .Y(N83) );
  NAND21X1 U42 ( .B(newinstr), .A(n9), .Y(n27) );
  OAI22X1 U43 ( .A(n8), .B(n31), .C(n59), .D(n27), .Y(n56) );
  NAND2X1 U44 ( .A(n12), .B(n26), .Y(t1ov) );
  NOR2X1 U45 ( .A(n31), .B(n14), .Y(n47) );
  NAND2X1 U46 ( .A(n38), .B(n9), .Y(n36) );
  NOR2X1 U47 ( .A(n8), .B(n38), .Y(N100) );
  AO22AXL U48 ( .A(n18), .B(n19), .C(t1_tf1), .D(n18), .Y(n54) );
  OAI31XL U49 ( .A(n20), .B(n8), .C(n7), .D(n21), .Y(n19) );
  OAI211X1 U50 ( .C(n22), .D(n21), .A(n20), .B(n23), .Y(n18) );
  NAND3X1 U51 ( .A(n24), .B(n20), .C(n23), .Y(n21) );
  AO222X1 U52 ( .A(n43), .B(th1[2]), .C(N44), .D(n44), .E(n45), .F(sfrdatai[2]), .Y(N53) );
  AO222X1 U53 ( .A(n43), .B(th1[3]), .C(N45), .D(n44), .E(n45), .F(sfrdatai[3]), .Y(N54) );
  AO222X1 U54 ( .A(n43), .B(th1[7]), .C(N49), .D(n44), .E(n45), .F(sfrdatai[7]), .Y(N58) );
  AO222X1 U55 ( .A(n43), .B(th1[6]), .C(N48), .D(n44), .E(n45), .F(sfrdatai[6]), .Y(N57) );
  AO222X1 U56 ( .A(n43), .B(th1[5]), .C(N47), .D(n44), .E(n45), .F(sfrdatai[5]), .Y(N56) );
  AO222X1 U57 ( .A(n43), .B(th1[4]), .C(N46), .D(n44), .E(n45), .F(sfrdatai[4]), .Y(N55) );
  AO222X1 U58 ( .A(n43), .B(th1[1]), .C(N43), .D(n44), .E(n45), .F(sfrdatai[1]), .Y(N52) );
  AO222X1 U59 ( .A(n43), .B(th1[0]), .C(N42), .D(n44), .E(n45), .F(sfrdatai[0]), .Y(N51) );
  ENOX1 U60 ( .A(n39), .B(n2), .C(N68), .D(n11), .Y(N77) );
  ENOX1 U61 ( .A(n7), .B(n39), .C(N75), .D(n11), .Y(N84) );
  NOR2X1 U62 ( .A(n8), .B(n32), .Y(n58) );
  AOI22AXL U63 ( .A(t1_tr1), .B(n20), .D(n20), .C(sfrdatai[6]), .Y(n32) );
  AO22AXL U64 ( .A(t1ack), .B(n9), .C(t1clr), .D(n27), .Y(n57) );
  OAI22AX1 U65 ( .D(th1_ov_ff), .C(n27), .A(n8), .B(n26), .Y(n55) );
  OAI2B11X1 U66 ( .D(t1_tmod[3]), .C(int1ff), .A(clk_ov12), .B(n51), .Y(n48)
         );
  AOI221XL U67 ( .A(n13), .B(n24), .C(t1_tmod[1]), .D(t1_tmod[0]), .E(
        t1_tmod[2]), .Y(n51) );
  INVX1 U68 ( .A(t1_tr1), .Y(n13) );
  NAND4X1 U69 ( .A(tl1[3]), .B(tl1[2]), .C(tl1[4]), .D(n49), .Y(n31) );
  NOR42XL U70 ( .C(tl1[1]), .D(tl1[0]), .A(n48), .B(n50), .Y(n49) );
  AOI32X1 U71 ( .A(tl1[6]), .B(tl1[5]), .C(tl1[7]), .D(n15), .E(n14), .Y(n50)
         );
  INVX1 U72 ( .A(t1_tmod[0]), .Y(n15) );
  AOI211X1 U73 ( .C(th1_ov_ff), .D(n14), .A(t1ov), .B(n25), .Y(n22) );
  NOR3XL U74 ( .A(n59), .B(t1_tmod[0]), .C(n14), .Y(n25) );
  NAND4X1 U75 ( .A(th1[3]), .B(th1[2]), .C(n28), .D(n29), .Y(n26) );
  AND4X1 U76 ( .A(th1[4]), .B(th1[5]), .C(th1[6]), .D(th1[7]), .Y(n29) );
  AND3X1 U77 ( .A(th1[1]), .B(n30), .C(th1[0]), .Y(n28) );
  NOR2X1 U78 ( .A(n31), .B(t1_tmod[1]), .Y(n30) );
  NAND2X1 U79 ( .A(t0_mode[1]), .B(t0_mode[0]), .Y(n24) );
  INVX1 U80 ( .A(t1_tmod[1]), .Y(n14) );
  NAND31X1 U81 ( .C(n36), .A(clk_count[1]), .B(clk_count[0]), .Y(n34) );
  AOI21BBXL U82 ( .B(clk_count[1]), .C(n36), .A(N95), .Y(n35) );
  OAI32X1 U83 ( .A(n16), .B(clk_count[3]), .C(n34), .D(n35), .E(n17), .Y(N98)
         );
  INVX1 U84 ( .A(clk_count[3]), .Y(n17) );
  NOR2X1 U85 ( .A(n36), .B(clk_count[0]), .Y(N95) );
  NOR3XL U86 ( .A(rst), .B(t1clr), .C(t1ack), .Y(n23) );
  OAI22X1 U87 ( .A(n35), .B(n16), .C(clk_count[2]), .D(n34), .Y(N97) );
  NOR2X1 U88 ( .A(n37), .B(n36), .Y(N96) );
  XNOR2XL U89 ( .A(clk_count[1]), .B(clk_count[0]), .Y(n37) );
  INVX1 U90 ( .A(tl1_ov_ff), .Y(n59) );
  NAND4X1 U91 ( .A(clk_count[3]), .B(clk_count[1]), .C(clk_count[0]), .D(n16), 
        .Y(n38) );
  INVX1 U92 ( .A(clk_count[2]), .Y(n16) );
endmodule


module timer1_a0_DW01_inc_1 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  XOR2X1 U1 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module timer1_a0_DW01_inc_0 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  XOR2X1 U1 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_timer1_a0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_timer1_a0_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_timer1_a0_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module timer0_a0 ( clkper, rst, newinstr, t0ff, t0ack, t1ack, int0ff, t0_tf0, 
        t0_tf1, sfrdatai, sfraddr, sfrwe, t0_tmod, t0_tr0, t0_tr1, tl0, th0 );
  input [7:0] sfrdatai;
  input [6:0] sfraddr;
  output [3:0] t0_tmod;
  output [7:0] tl0;
  output [7:0] th0;
  input clkper, rst, newinstr, t0ff, t0ack, t1ack, int0ff, sfrwe;
  output t0_tf0, t0_tf1, t0_tr0, t0_tr1;
  wire   t0clr, th0_ov_ff, tl0_ov_ff, t1clr, N39, N40, N41, N42, N43, N47, N48,
         N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62,
         N63, N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83,
         N84, N85, N86, N87, N101, N102, N103, N104, clk_ov12, N106, net12221,
         net12227, net12232, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n1, n2, n3, n4, n5, n6,
         n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n68, n69;
  wire   [3:0] clk_count;

  SNPS_CLOCK_GATE_HIGH_timer0_a0_0 clk_gate_t0_ct_reg ( .CLK(clkper), .EN(N39), 
        .ENCLK(net12221), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_timer0_a0_2 clk_gate_th0_s_reg ( .CLK(clkper), .EN(N55), 
        .ENCLK(net12227), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_timer0_a0_1 clk_gate_tl0_s_reg ( .CLK(clkper), .EN(N79), 
        .ENCLK(net12232), .TE(1'b0) );
  timer0_a0_DW01_inc_0 add_347 ( .A(tl0), .SUM({N78, N77, N76, N75, N74, N73, 
        N72, N71}) );
  timer0_a0_DW01_inc_1 add_309 ( .A(th0), .SUM({N54, N53, N52, N51, N50, N49, 
        N48, N47}) );
  DFFQX1 t1clr_reg ( .D(n63), .C(clkper), .Q(t1clr) );
  DFFQX1 clk_count_reg_1_ ( .D(N102), .C(clkper), .Q(clk_count[1]) );
  DFFQX1 tl0_ov_ff_reg ( .D(n64), .C(clkper), .Q(tl0_ov_ff) );
  DFFQX1 th0_ov_ff_reg ( .D(n61), .C(clkper), .Q(th0_ov_ff) );
  DFFQX1 clk_count_reg_2_ ( .D(N103), .C(clkper), .Q(clk_count[2]) );
  DFFQX1 clk_count_reg_0_ ( .D(N101), .C(clkper), .Q(clk_count[0]) );
  DFFQX1 t0clr_reg ( .D(n65), .C(clkper), .Q(t0clr) );
  DFFQX1 clk_count_reg_3_ ( .D(N104), .C(clkper), .Q(clk_count[3]) );
  DFFQX1 clk_ov12_reg ( .D(N106), .C(clkper), .Q(clk_ov12) );
  DFFQX1 tl0_s_reg_7_ ( .D(N87), .C(net12232), .Q(tl0[7]) );
  DFFQX1 tl0_s_reg_1_ ( .D(N81), .C(net12232), .Q(tl0[1]) );
  DFFQX1 t0_gate_reg ( .D(N40), .C(net12221), .Q(t0_tmod[3]) );
  DFFQX1 tl0_s_reg_3_ ( .D(N83), .C(net12232), .Q(tl0[3]) );
  DFFQX1 t0_tf0_s_reg ( .D(n60), .C(clkper), .Q(t0_tf0) );
  DFFQX1 th0_s_reg_2_ ( .D(N58), .C(net12227), .Q(th0[2]) );
  DFFQX1 t0_ct_reg ( .D(N41), .C(net12221), .Q(t0_tmod[2]) );
  DFFQX1 tl0_s_reg_2_ ( .D(N82), .C(net12232), .Q(tl0[2]) );
  DFFQX1 t0_mode_reg_1_ ( .D(N43), .C(net12221), .Q(t0_tmod[1]) );
  DFFQX1 t0_tf1_s_reg ( .D(n62), .C(clkper), .Q(t0_tf1) );
  DFFQX1 t0_tr1_s_reg ( .D(n66), .C(clkper), .Q(t0_tr1) );
  DFFQX1 tl0_s_reg_5_ ( .D(N85), .C(net12232), .Q(tl0[5]) );
  DFFQX1 tl0_s_reg_6_ ( .D(N86), .C(net12232), .Q(tl0[6]) );
  DFFQX1 tl0_s_reg_0_ ( .D(N80), .C(net12232), .Q(tl0[0]) );
  DFFQX1 th0_s_reg_7_ ( .D(N63), .C(net12227), .Q(th0[7]) );
  DFFQX1 t0_tr0_s_reg ( .D(n67), .C(clkper), .Q(t0_tr0) );
  DFFQX1 th0_s_reg_5_ ( .D(N61), .C(net12227), .Q(th0[5]) );
  DFFQX1 th0_s_reg_4_ ( .D(N60), .C(net12227), .Q(th0[4]) );
  DFFQX1 th0_s_reg_6_ ( .D(N62), .C(net12227), .Q(th0[6]) );
  DFFQX1 th0_s_reg_1_ ( .D(N57), .C(net12227), .Q(th0[1]) );
  DFFQX1 tl0_s_reg_4_ ( .D(N84), .C(net12232), .Q(tl0[4]) );
  DFFQX1 th0_s_reg_0_ ( .D(N56), .C(net12227), .Q(th0[0]) );
  DFFQX1 th0_s_reg_3_ ( .D(N59), .C(net12227), .Q(th0[3]) );
  DFFQX1 t0_mode_reg_0_ ( .D(N42), .C(net12221), .Q(t0_tmod[0]) );
  NOR2X1 U3 ( .A(n11), .B(n34), .Y(n23) );
  NAND21X1 U4 ( .B(n48), .A(n10), .Y(n47) );
  INVX1 U5 ( .A(n34), .Y(n13) );
  NAND2X1 U6 ( .A(n10), .B(n53), .Y(N39) );
  INVX1 U7 ( .A(rst), .Y(n10) );
  NOR21XL U8 ( .B(n52), .A(sfraddr[2]), .Y(n39) );
  NOR2X1 U9 ( .A(n26), .B(n11), .Y(n34) );
  NAND3X1 U10 ( .A(n1), .B(n2), .C(n39), .Y(n26) );
  NOR2X1 U11 ( .A(n45), .B(n11), .Y(n42) );
  NAND4X1 U12 ( .A(sfraddr[2]), .B(n52), .C(n1), .D(n2), .Y(n48) );
  NAND4X1 U13 ( .A(sfraddr[0]), .B(n39), .C(n10), .D(n2), .Y(n53) );
  NOR2X1 U14 ( .A(n6), .B(n53), .Y(N40) );
  NOR2X1 U15 ( .A(n3), .B(n53), .Y(N42) );
  NOR2X1 U16 ( .A(n4), .B(n53), .Y(N43) );
  NOR2X1 U17 ( .A(n5), .B(n53), .Y(N41) );
  INVX1 U18 ( .A(sfraddr[0]), .Y(n1) );
  INVX1 U19 ( .A(n12), .Y(n11) );
  AND3X1 U20 ( .A(sfrwe), .B(sfraddr[3]), .C(n54), .Y(n52) );
  NOR3XL U21 ( .A(sfraddr[4]), .B(sfraddr[6]), .C(sfraddr[5]), .Y(n54) );
  OR4X1 U22 ( .A(n42), .B(n40), .C(n41), .D(n11), .Y(N79) );
  NAND3X1 U23 ( .A(n39), .B(n1), .C(sfraddr[1]), .Y(n45) );
  NAND32X1 U24 ( .B(n46), .C(n11), .A(n47), .Y(N55) );
  INVX1 U25 ( .A(sfraddr[1]), .Y(n2) );
  INVX1 U26 ( .A(sfrdatai[3]), .Y(n6) );
  INVX1 U27 ( .A(sfrdatai[0]), .Y(n3) );
  INVX1 U28 ( .A(sfrdatai[1]), .Y(n4) );
  INVX1 U29 ( .A(sfrdatai[2]), .Y(n5) );
  INVX1 U30 ( .A(sfrdatai[6]), .Y(n9) );
  INVX1 U31 ( .A(sfrdatai[4]), .Y(n7) );
  INVX1 U32 ( .A(sfrdatai[5]), .Y(n8) );
  INVX1 U33 ( .A(rst), .Y(n12) );
  INVX1 U34 ( .A(t0ack), .Y(n14) );
  NOR32XL U35 ( .B(n45), .C(n10), .A(n44), .Y(n40) );
  AND4X1 U36 ( .A(n43), .B(n44), .C(n45), .D(n10), .Y(n41) );
  NOR32XL U37 ( .B(n48), .C(n10), .A(n38), .Y(n46) );
  ENOX1 U38 ( .A(n9), .B(n47), .C(N53), .D(n46), .Y(N62) );
  ENOX1 U39 ( .A(n8), .B(n47), .C(N52), .D(n46), .Y(N61) );
  ENOX1 U40 ( .A(n7), .B(n47), .C(N51), .D(n46), .Y(N60) );
  ENOX1 U41 ( .A(n6), .B(n47), .C(N50), .D(n46), .Y(N59) );
  ENOX1 U42 ( .A(n5), .B(n47), .C(N49), .D(n46), .Y(N58) );
  ENOX1 U43 ( .A(n4), .B(n47), .C(N48), .D(n46), .Y(N57) );
  NAND21X1 U44 ( .B(newinstr), .A(n10), .Y(n30) );
  OAI22X1 U45 ( .A(n11), .B(n14), .C(n30), .D(n20), .Y(n65) );
  OAI22X1 U46 ( .A(n11), .B(n29), .C(n30), .D(n69), .Y(n61) );
  OAI22X1 U47 ( .A(n11), .B(n28), .C(n30), .D(n68), .Y(n64) );
  INVX1 U48 ( .A(n28), .Y(n15) );
  NAND2X1 U49 ( .A(n55), .B(n10), .Y(n58) );
  NOR2X1 U50 ( .A(n16), .B(n17), .Y(n35) );
  NOR2X1 U51 ( .A(n11), .B(n55), .Y(N106) );
  OAI22BX1 U52 ( .B(n31), .A(n32), .D(t0_tf1), .C(n31), .Y(n62) );
  AOI32X1 U53 ( .A(n26), .B(n10), .C(n33), .D(sfrdatai[7]), .E(n34), .Y(n32)
         );
  OAI2B11X1 U54 ( .D(n35), .C(n29), .A(n23), .B(n33), .Y(n31) );
  NOR2X1 U55 ( .A(t1clr), .B(t1ack), .Y(n33) );
  OAI211X1 U56 ( .C(n13), .D(n8), .A(n21), .B(n22), .Y(n60) );
  OAI211X1 U57 ( .C(n24), .D(n25), .A(n26), .B(n27), .Y(n21) );
  NAND4X1 U58 ( .A(t0_tf0), .B(n23), .C(n14), .D(n20), .Y(n22) );
  AOI21X1 U59 ( .B(n68), .C(n28), .A(n16), .Y(n25) );
  AO222X1 U60 ( .A(n40), .B(th0[7]), .C(N78), .D(n41), .E(n42), .F(sfrdatai[7]), .Y(N87) );
  AO222X1 U61 ( .A(n40), .B(th0[6]), .C(N77), .D(n41), .E(n42), .F(sfrdatai[6]), .Y(N86) );
  AO222X1 U62 ( .A(n40), .B(th0[5]), .C(N76), .D(n41), .E(n42), .F(sfrdatai[5]), .Y(N85) );
  AO222X1 U63 ( .A(n40), .B(th0[4]), .C(N75), .D(n41), .E(n42), .F(sfrdatai[4]), .Y(N84) );
  AO222X1 U64 ( .A(n40), .B(th0[3]), .C(N74), .D(n41), .E(sfrdatai[3]), .F(n42), .Y(N83) );
  AO222X1 U65 ( .A(n40), .B(th0[2]), .C(N73), .D(n41), .E(sfrdatai[2]), .F(n42), .Y(N82) );
  AO222X1 U66 ( .A(n40), .B(th0[1]), .C(N72), .D(n41), .E(sfrdatai[1]), .F(n42), .Y(N81) );
  AO222X1 U67 ( .A(n40), .B(th0[0]), .C(N71), .D(n41), .E(sfrdatai[0]), .F(n42), .Y(N80) );
  AO22AXL U68 ( .A(N54), .B(n46), .C(sfrdatai[7]), .D(n47), .Y(N63) );
  ENOX1 U69 ( .A(n13), .B(n9), .C(t0_tr1), .D(n23), .Y(n66) );
  ENOX1 U70 ( .A(n13), .B(n7), .C(t0_tr0), .D(n23), .Y(n67) );
  ENOX1 U71 ( .A(n3), .B(n47), .C(N47), .D(n46), .Y(N56) );
  AO22AXL U72 ( .A(t1ack), .B(n10), .C(t1clr), .D(n30), .Y(n63) );
  NAND4X1 U73 ( .A(tl0[3]), .B(tl0[2]), .C(tl0[4]), .D(n49), .Y(n28) );
  NOR43XL U74 ( .B(tl0[1]), .C(tl0[0]), .D(n43), .A(n50), .Y(n49) );
  AOI32X1 U75 ( .A(tl0[6]), .B(tl0[5]), .C(tl0[7]), .D(n17), .E(n16), .Y(n50)
         );
  NOR43XL U76 ( .B(clk_ov12), .C(n51), .D(t0_tr0), .A(t0_tmod[2]), .Y(n43) );
  NAND21X1 U77 ( .B(int0ff), .A(t0_tmod[3]), .Y(n51) );
  AOI32X1 U78 ( .A(t0_tr1), .B(n35), .C(clk_ov12), .D(n16), .E(n15), .Y(n38)
         );
  INVX1 U79 ( .A(t0_tmod[1]), .Y(n16) );
  AOI21X1 U80 ( .B(n69), .C(n29), .A(t0_tmod[1]), .Y(n24) );
  NAND4X1 U81 ( .A(th0[3]), .B(th0[2]), .C(n36), .D(n37), .Y(n29) );
  AND4X1 U82 ( .A(th0[4]), .B(th0[5]), .C(th0[6]), .D(th0[7]), .Y(n37) );
  NOR32XL U83 ( .B(th0[1]), .C(th0[0]), .A(n38), .Y(n36) );
  INVX1 U84 ( .A(t0_tmod[0]), .Y(n17) );
  NAND31X1 U85 ( .C(n58), .A(clk_count[1]), .B(clk_count[0]), .Y(n56) );
  AOI21BBXL U86 ( .B(clk_count[1]), .C(n58), .A(N101), .Y(n57) );
  OAI32X1 U87 ( .A(n18), .B(clk_count[3]), .C(n56), .D(n57), .E(n19), .Y(N104)
         );
  INVX1 U88 ( .A(clk_count[3]), .Y(n19) );
  NOR2X1 U89 ( .A(n58), .B(clk_count[0]), .Y(N101) );
  OAI22X1 U90 ( .A(n57), .B(n18), .C(clk_count[2]), .D(n56), .Y(N103) );
  NAND3X1 U91 ( .A(t0_tmod[1]), .B(n17), .C(n15), .Y(n44) );
  NOR3XL U92 ( .A(n11), .B(t0clr), .C(t0ack), .Y(n27) );
  NOR2X1 U93 ( .A(n59), .B(n58), .Y(N102) );
  XNOR2XL U94 ( .A(clk_count[1]), .B(clk_count[0]), .Y(n59) );
  NAND4X1 U95 ( .A(clk_count[3]), .B(clk_count[1]), .C(clk_count[0]), .D(n18), 
        .Y(n55) );
  INVX1 U96 ( .A(clk_count[2]), .Y(n18) );
  INVX1 U97 ( .A(th0_ov_ff), .Y(n69) );
  INVX1 U98 ( .A(tl0_ov_ff), .Y(n68) );
  INVX1 U99 ( .A(t0clr), .Y(n20) );
endmodule


module timer0_a0_DW01_inc_1 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  XOR2X1 U1 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module timer0_a0_DW01_inc_0 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  XOR2X1 U1 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_timer0_a0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_timer0_a0_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_timer0_a0_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module serial0_a0 ( t_shift_clk, r_shift_clk, clkper, rst, newinstr, rxd0ff, 
        t1ov, rxd0o, rxd0oe, txd0, sfrdatai, sfraddr, sfrwe, s0con, s0buf, 
        s0rell, s0relh, smod, bd );
  input [7:0] sfrdatai;
  input [6:0] sfraddr;
  output [7:0] s0con;
  output [7:0] s0buf;
  output [7:0] s0rell;
  output [7:0] s0relh;
  input clkper, rst, newinstr, rxd0ff, t1ov, sfrwe;
  output t_shift_clk, r_shift_clk, rxd0o, rxd0oe, txd0, smod, bd;
  wire   r_clk_ov2, t1ov_ff, N59, ri_tmp, rxd0_val, s0con2_val, s0con2_tmp,
         ti_tmp, N108, N109, N110, N111, N112, N113, N117, N118, N119, N120,
         N121, N122, N123, N124, N125, N128, N129, N130, N131, N132, N133,
         N134, N135, N136, baud_rate_ov, N142, N145, N146, N147, N148, N149,
         N150, N151, N152, N153, N154, N166, N169, N170, N185, N186, N187,
         N188, N190, clk_ov12, N191, r_start, baud_r_count, baud_r2_clk, N207,
         t_baud_ov, t_start, N223, N224, N225, N226, N227, N230, N257, N258,
         N259, N260, N261, N262, N263, N264, N265, N266, N267, N268, N281,
         N282, N283, N284, N303, rxd0_fall, rxd0_ff, rxd0_fall_fl,
         receive_11_bits, N306, N307, N324, N325, N326, N327, N333, ri0_fall,
         ri0_ff, N348, N360, N361, N362, N363, N364, N375, N376, N377, N378,
         N379, N380, N381, N382, N424, N425, N426, N427, N428, N471, N472,
         N473, N474, N475, N476, N477, N478, N479, net12260, net12266,
         net12271, net12276, net12281, net12286, net12291, net12296, net12301,
         net12306, net12311, n13, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n1, n2, n3, n4, n5, n6, n7, n8,
         n9, n10, n11, n12, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256;
  wire   [3:0] r_baud_count;
  wire   [3:0] r_shift_count;
  wire   [3:0] t_shift_count;
  wire   [9:0] tim_baud;
  wire   [3:0] clk_count;
  wire   [3:0] t_baud_count;
  wire   [10:0] t_shift_reg;
  wire   [1:0] fluctuation_conter;
  wire   [2:0] rxd0_vec;
  wire   [7:0] r_shift_reg;

  MAJ3X1 U336 ( .A(rxd0_vec[1]), .B(rxd0_vec[0]), .C(rxd0_vec[2]), .Y(n172) );
  SNPS_CLOCK_GATE_HIGH_serial0_a0_0 clk_gate_s0con_s_reg ( .CLK(clkper), .EN(
        N108), .ENCLK(net12260), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_serial0_a0_10 clk_gate_s0rell_s_reg ( .CLK(clkper), 
        .EN(N117), .ENCLK(net12266), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_serial0_a0_9 clk_gate_s0relh_s_reg ( .CLK(clkper), .EN(
        N128), .ENCLK(net12271), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_serial0_a0_8 clk_gate_tim_baud_reg ( .CLK(clkper), .EN(
        N166), .ENCLK(net12276), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_serial0_a0_7 clk_gate_t_baud_count_reg ( .CLK(clkper), 
        .EN(N223), .ENCLK(net12281), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_serial0_a0_6 clk_gate_t_shift_reg_reg ( .CLK(clkper), 
        .EN(N257), .ENCLK(net12286), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_serial0_a0_5 clk_gate_rxd0_vec_reg ( .CLK(clkper), .EN(
        N324), .ENCLK(net12291), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_serial0_a0_4 clk_gate_r_baud_count_reg ( .CLK(clkper), 
        .EN(N360), .ENCLK(net12296), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_serial0_a0_3 clk_gate_r_shift_reg_reg ( .CLK(clkper), 
        .EN(n13), .ENCLK(net12301), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_serial0_a0_2 clk_gate_r_shift_count_reg ( .CLK(clkper), 
        .EN(N428), .ENCLK(net12306), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_serial0_a0_1 clk_gate_s0buf_r_reg ( .CLK(clkper), .EN(
        N471), .ENCLK(net12311), .TE(1'b0) );
  serial0_a0_DW01_inc_0 add_584 ( .A(tim_baud), .SUM({N154, N153, N152, N151, 
        N150, N149, N148, N147, N146, N145}) );
  DFFQX1 t_shift_reg_reg_9_ ( .D(N267), .C(net12286), .Q(t_shift_reg[9]) );
  DFFQX1 t_shift_reg_reg_8_ ( .D(N266), .C(net12286), .Q(t_shift_reg[8]) );
  DFFQX1 t_shift_reg_reg_7_ ( .D(N265), .C(net12286), .Q(t_shift_reg[7]) );
  DFFQX1 t_shift_reg_reg_6_ ( .D(N264), .C(net12286), .Q(t_shift_reg[6]) );
  DFFQX1 t_shift_reg_reg_5_ ( .D(N263), .C(net12286), .Q(t_shift_reg[5]) );
  DFFQX1 t_shift_reg_reg_4_ ( .D(N262), .C(net12286), .Q(t_shift_reg[4]) );
  DFFQX1 t_shift_reg_reg_3_ ( .D(N261), .C(net12286), .Q(t_shift_reg[3]) );
  DFFQX1 t_shift_reg_reg_10_ ( .D(N268), .C(net12286), .Q(t_shift_reg[10]) );
  DFFQX1 r_shift_reg_reg_0_ ( .D(N375), .C(net12301), .Q(r_shift_reg[0]) );
  DFFQX1 t_shift_reg_reg_1_ ( .D(N259), .C(net12286), .Q(t_shift_reg[1]) );
  DFFQX1 rxd0_vec_reg_2_ ( .D(N327), .C(net12291), .Q(rxd0_vec[2]) );
  DFFQX1 rxd0_vec_reg_1_ ( .D(N326), .C(net12291), .Q(rxd0_vec[1]) );
  DFFQX1 t_shift_reg_reg_0_ ( .D(N258), .C(net12286), .Q(t_shift_reg[0]) );
  DFFQX1 ti_tmp_reg ( .D(n242), .C(clkper), .Q(ti_tmp) );
  DFFQX1 rxd0_ff_reg ( .D(N307), .C(clkper), .Q(rxd0_ff) );
  DFFQX1 t_shift_reg_reg_2_ ( .D(N260), .C(net12286), .Q(t_shift_reg[2]) );
  DFFQX1 rxd0_vec_reg_0_ ( .D(N325), .C(net12291), .Q(rxd0_vec[0]) );
  DFFQX1 baud_r_count_reg ( .D(n245), .C(clkper), .Q(baud_r_count) );
  DFFQX1 r_shift_reg_reg_7_ ( .D(N382), .C(net12301), .Q(r_shift_reg[7]) );
  DFFQX1 r_shift_reg_reg_6_ ( .D(N381), .C(net12301), .Q(r_shift_reg[6]) );
  DFFQX1 r_shift_reg_reg_5_ ( .D(N380), .C(net12301), .Q(r_shift_reg[5]) );
  DFFQX1 r_shift_reg_reg_4_ ( .D(N379), .C(net12301), .Q(r_shift_reg[4]) );
  DFFQX1 r_shift_reg_reg_3_ ( .D(N378), .C(net12301), .Q(r_shift_reg[3]) );
  DFFQX1 r_shift_reg_reg_2_ ( .D(N377), .C(net12301), .Q(r_shift_reg[2]) );
  DFFQX1 r_shift_reg_reg_1_ ( .D(N376), .C(net12301), .Q(r_shift_reg[1]) );
  DFFQX1 ri_tmp_reg ( .D(n238), .C(clkper), .Q(ri_tmp) );
  DFFQX1 fluctuation_conter_reg_0_ ( .D(n234), .C(clkper), .Q(
        fluctuation_conter[0]) );
  DFFQX1 s0con2_val_reg ( .D(n231), .C(net12291), .Q(s0con2_val) );
  DFFQX1 s0con2_tmp_reg ( .D(n232), .C(clkper), .Q(s0con2_tmp) );
  DFFQX1 receive_11_bits_reg ( .D(n229), .C(clkper), .Q(receive_11_bits) );
  DFFQX1 fluctuation_conter_reg_1_ ( .D(n233), .C(clkper), .Q(
        fluctuation_conter[1]) );
  DFFQX1 ri0_fall_reg ( .D(n236), .C(clkper), .Q(ri0_fall) );
  DFFQX1 ri0_ff_reg ( .D(N348), .C(clkper), .Q(ri0_ff) );
  DFFQX1 t_shift_count_reg_1_ ( .D(N282), .C(net12286), .Q(t_shift_count[1])
         );
  DFFQX1 rxd0_fall_fl_reg ( .D(n235), .C(clkper), .Q(rxd0_fall_fl) );
  DFFQX1 t_shift_count_reg_3_ ( .D(N284), .C(net12286), .Q(t_shift_count[3])
         );
  DFFQX1 t_shift_count_reg_2_ ( .D(N283), .C(net12286), .Q(t_shift_count[2])
         );
  DFFQX1 clk_count_reg_1_ ( .D(N186), .C(clkper), .Q(clk_count[1]) );
  DFFQX1 t_shift_count_reg_0_ ( .D(N281), .C(net12286), .Q(t_shift_count[0])
         );
  DFFQX1 clk_count_reg_0_ ( .D(N185), .C(clkper), .Q(clk_count[0]) );
  DFFQX1 rxd0_val_reg ( .D(N333), .C(clkper), .Q(rxd0_val) );
  DFFQX1 clk_count_reg_3_ ( .D(N188), .C(clkper), .Q(clk_count[3]) );
  DFFQX1 clk_count_reg_2_ ( .D(N187), .C(clkper), .Q(clk_count[2]) );
  DFFQX1 rxd0_fall_reg ( .D(N306), .C(clkper), .Q(rxd0_fall) );
  DFFQX1 clk_ov12_reg ( .D(N191), .C(clkper), .Q(clk_ov12) );
  DFFQX1 t_baud_ov_reg ( .D(N230), .C(clkper), .Q(t_baud_ov) );
  DFFQX1 baud_r2_clk_reg ( .D(N207), .C(clkper), .Q(baud_r2_clk) );
  DFFQX1 tim_baud_reg_9_ ( .D(n62), .C(net12276), .Q(tim_baud[9]) );
  DFFQX1 tim_baud_reg_8_ ( .D(n61), .C(net12276), .Q(tim_baud[8]) );
  DFFQX1 tim_baud_reg_3_ ( .D(N170), .C(net12276), .Q(tim_baud[3]) );
  DFFQX1 tim_baud_reg_4_ ( .D(n58), .C(net12276), .Q(tim_baud[4]) );
  DFFQX1 t_baud_count_reg_3_ ( .D(N227), .C(net12281), .Q(t_baud_count[3]) );
  DFFQX1 r_baud_count_reg_3_ ( .D(N364), .C(net12296), .Q(r_baud_count[3]) );
  DFFQX1 r_shift_count_reg_1_ ( .D(N425), .C(net12306), .Q(r_shift_count[1])
         );
  DFFQX1 r_shift_count_reg_3_ ( .D(N427), .C(net12306), .Q(r_shift_count[3])
         );
  DFFQX1 r_shift_count_reg_2_ ( .D(N426), .C(net12306), .Q(r_shift_count[2])
         );
  DFFQX1 t_baud_count_reg_1_ ( .D(N225), .C(net12281), .Q(t_baud_count[1]) );
  DFFQX1 t_baud_count_reg_0_ ( .D(N224), .C(net12281), .Q(t_baud_count[0]) );
  DFFQX1 t_baud_count_reg_2_ ( .D(N226), .C(net12281), .Q(t_baud_count[2]) );
  DFFQX1 r_start_reg ( .D(n240), .C(clkper), .Q(r_start) );
  DFFQX1 t1ov_ff_reg ( .D(N59), .C(clkper), .Q(t1ov_ff) );
  DFFQX1 tim_baud_reg_2_ ( .D(N169), .C(net12276), .Q(tim_baud[2]) );
  DFFQX1 tim_baud_reg_7_ ( .D(n55), .C(net12276), .Q(tim_baud[7]) );
  DFFQX1 tim_baud_reg_5_ ( .D(n57), .C(net12276), .Q(tim_baud[5]) );
  DFFQX1 tim_baud_reg_1_ ( .D(n59), .C(net12276), .Q(tim_baud[1]) );
  DFFQX1 tim_baud_reg_6_ ( .D(n56), .C(net12276), .Q(tim_baud[6]) );
  DFFQX1 tim_baud_reg_0_ ( .D(n60), .C(net12276), .Q(tim_baud[0]) );
  DFFQX1 r_baud_count_reg_1_ ( .D(N362), .C(net12296), .Q(r_baud_count[1]) );
  DFFQX1 r_shift_count_reg_0_ ( .D(N424), .C(net12306), .Q(r_shift_count[0])
         );
  DFFQX1 r_baud_count_reg_2_ ( .D(N363), .C(net12296), .Q(r_baud_count[2]) );
  DFFQX1 r_baud_count_reg_0_ ( .D(N361), .C(net12296), .Q(r_baud_count[0]) );
  DFFQX1 baud_rate_ov_reg ( .D(N142), .C(clkper), .Q(baud_rate_ov) );
  DFFQX1 r_clk_ov2_reg ( .D(N190), .C(clkper), .Q(r_clk_ov2) );
  DFFQX1 rxd0o_reg ( .D(N303), .C(clkper), .Q(rxd0o) );
  DFFQX1 t_start_reg ( .D(n243), .C(clkper), .Q(t_start) );
  DFFQX1 txd0_reg ( .D(n239), .C(clkper), .Q(txd0) );
  DFFQX1 s0relh_s_reg_5_ ( .D(N134), .C(net12271), .Q(s0relh[5]) );
  DFFQX1 s0relh_s_reg_4_ ( .D(N133), .C(net12271), .Q(s0relh[4]) );
  DFFQX1 s0relh_s_reg_3_ ( .D(N132), .C(net12271), .Q(s0relh[3]) );
  DFFQX1 s0buf_r_reg_7_ ( .D(N479), .C(net12311), .Q(s0buf[7]) );
  DFFQX1 s0buf_r_reg_2_ ( .D(N474), .C(net12311), .Q(s0buf[2]) );
  DFFQX1 s0rell_s_reg_2_ ( .D(N120), .C(net12266), .Q(s0rell[2]) );
  DFFQX1 s0rell_s_reg_3_ ( .D(N121), .C(net12266), .Q(s0rell[3]) );
  DFFQX1 s0relh_s_reg_1_ ( .D(N130), .C(net12271), .Q(s0relh[1]) );
  DFFQX1 s0relh_s_reg_0_ ( .D(N129), .C(net12271), .Q(s0relh[0]) );
  DFFQX1 s0rell_s_reg_1_ ( .D(N119), .C(net12266), .Q(s0rell[1]) );
  DFFQX1 s0rell_s_reg_7_ ( .D(N125), .C(net12266), .Q(s0rell[7]) );
  DFFQX1 s0relh_s_reg_2_ ( .D(N131), .C(net12271), .Q(s0relh[2]) );
  DFFQX1 bd_s_reg ( .D(n42), .C(clkper), .Q(bd) );
  DFFQX1 smod_s_reg ( .D(n244), .C(clkper), .Q(smod) );
  DFFQX1 s0con_s_reg_2_ ( .D(n230), .C(clkper), .Q(s0con[2]) );
  DFFQX1 s0relh_s_reg_7_ ( .D(N136), .C(net12271), .Q(s0relh[7]) );
  DFFQX1 s0relh_s_reg_6_ ( .D(N135), .C(net12271), .Q(s0relh[6]) );
  DFFQX1 s0buf_r_reg_5_ ( .D(N477), .C(net12311), .Q(s0buf[5]) );
  DFFQX1 s0buf_r_reg_4_ ( .D(N476), .C(net12311), .Q(s0buf[4]) );
  DFFQX1 s0buf_r_reg_0_ ( .D(N472), .C(net12311), .Q(s0buf[0]) );
  DFFQX1 s0buf_r_reg_6_ ( .D(N478), .C(net12311), .Q(s0buf[6]) );
  DFFQX1 s0buf_r_reg_3_ ( .D(N475), .C(net12311), .Q(s0buf[3]) );
  DFFQX1 s0buf_r_reg_1_ ( .D(N473), .C(net12311), .Q(s0buf[1]) );
  DFFQX1 s0con_s_reg_3_ ( .D(N109), .C(net12260), .Q(s0con[3]) );
  DFFQX1 s0rell_s_reg_5_ ( .D(N123), .C(net12266), .Q(s0rell[5]) );
  DFFQX1 s0rell_s_reg_4_ ( .D(N122), .C(net12266), .Q(s0rell[4]) );
  DFFQX1 s0rell_s_reg_0_ ( .D(N118), .C(net12266), .Q(s0rell[0]) );
  DFFQX1 s0con_s_reg_1_ ( .D(n241), .C(clkper), .Q(s0con[1]) );
  DFFQX1 s0con_s_reg_5_ ( .D(N111), .C(net12260), .Q(s0con[5]) );
  DFFQX1 s0con_s_reg_4_ ( .D(N110), .C(net12260), .Q(s0con[4]) );
  DFFQX1 s0con_s_reg_0_ ( .D(n237), .C(clkper), .Q(s0con[0]) );
  DFFQX1 s0con_s_reg_6_ ( .D(N112), .C(net12260), .Q(s0con[6]) );
  DFFQX1 s0con_s_reg_7_ ( .D(N113), .C(net12260), .Q(s0con[7]) );
  DFFQX1 s0rell_s_reg_6_ ( .D(N124), .C(net12266), .Q(s0rell[6]) );
  INVX1 U3 ( .A(n221), .Y(n1) );
  BUFX3 U4 ( .A(n211), .Y(n2) );
  INVX1 U5 ( .A(n51), .Y(n3) );
  NAND31XL U6 ( .C(sfraddr[6]), .A(n4), .B(n146), .Y(n134) );
  AOI221XL U7 ( .A(n87), .B(r_shift_clk), .C(r_start), .D(n49), .E(n28), .Y(
        n151) );
  AOI22AXL U8 ( .A(n64), .B(baud_rate_ov), .D(n222), .C(s0relh[7]), .Y(n221)
         );
  INVX1 U9 ( .A(N108), .Y(n39) );
  NAND2X1 U10 ( .A(n15), .B(n40), .Y(N108) );
  INVX1 U11 ( .A(n133), .Y(n40) );
  INVX1 U12 ( .A(n183), .Y(n36) );
  INVX1 U13 ( .A(n113), .Y(n41) );
  INVX1 U14 ( .A(n181), .Y(n35) );
  INVX1 U15 ( .A(n21), .Y(n15) );
  INVX1 U16 ( .A(n24), .Y(n16) );
  INVX1 U17 ( .A(n25), .Y(n17) );
  INVX1 U18 ( .A(n24), .Y(n18) );
  INVX1 U19 ( .A(n20), .Y(n19) );
  NOR2X1 U20 ( .A(n193), .B(n22), .Y(n181) );
  NOR2X1 U21 ( .A(n134), .B(n22), .Y(n133) );
  NOR4XL U22 ( .A(n44), .B(n5), .C(sfraddr[0]), .D(sfraddr[2]), .Y(n227) );
  NAND2X1 U23 ( .A(n181), .B(n51), .Y(n183) );
  NAND2X1 U24 ( .A(n134), .B(n15), .Y(n113) );
  INVX1 U25 ( .A(n176), .Y(n38) );
  OAI21X1 U26 ( .B(n40), .C(n12), .A(n19), .Y(N112) );
  OAI21X1 U27 ( .B(n6), .C(n226), .A(n19), .Y(N129) );
  OAI21X1 U28 ( .B(n7), .C(n226), .A(n19), .Y(N130) );
  OAI21X1 U29 ( .B(n6), .C(n228), .A(n19), .Y(N118) );
  OAI21X1 U30 ( .B(n9), .C(n228), .A(n19), .Y(N121) );
  OAI21X1 U31 ( .B(n10), .C(n228), .A(n19), .Y(N122) );
  OAI21X1 U32 ( .B(n12), .C(n228), .A(n31), .Y(N124) );
  OAI21X1 U33 ( .B(n14), .C(n228), .A(n31), .Y(N125) );
  NOR2X1 U34 ( .A(n7), .B(n228), .Y(N119) );
  NOR2X1 U35 ( .A(n8), .B(n228), .Y(N120) );
  NOR2X1 U36 ( .A(n11), .B(n228), .Y(N123) );
  NOR2X1 U37 ( .A(n8), .B(n226), .Y(N131) );
  NOR2X1 U38 ( .A(n9), .B(n226), .Y(N132) );
  NOR2X1 U39 ( .A(n10), .B(n226), .Y(N133) );
  NOR2X1 U40 ( .A(n11), .B(n226), .Y(N134) );
  NOR2X1 U41 ( .A(n12), .B(n226), .Y(N135) );
  NOR2X1 U42 ( .A(n14), .B(n226), .Y(N136) );
  NOR2X1 U43 ( .A(n40), .B(n9), .Y(N109) );
  NOR2X1 U44 ( .A(n40), .B(n10), .Y(N110) );
  NOR2X1 U45 ( .A(n40), .B(n11), .Y(N111) );
  NOR2X1 U46 ( .A(n40), .B(n14), .Y(N113) );
  NAND3X1 U47 ( .A(n35), .B(n17), .C(n176), .Y(N257) );
  NAND2X1 U48 ( .A(n16), .B(n226), .Y(N128) );
  NAND2X1 U49 ( .A(n15), .B(n228), .Y(N117) );
  INVX1 U50 ( .A(n30), .Y(n24) );
  INVX1 U51 ( .A(n31), .Y(n21) );
  INVX1 U52 ( .A(n30), .Y(n25) );
  INVX1 U53 ( .A(n29), .Y(n22) );
  INVX1 U54 ( .A(n19), .Y(n23) );
  INVX1 U55 ( .A(n29), .Y(n26) );
  INVX1 U56 ( .A(n29), .Y(n27) );
  INVX1 U57 ( .A(n31), .Y(n20) );
  INVX1 U58 ( .A(n29), .Y(n28) );
  INVX1 U59 ( .A(n112), .Y(n49) );
  INVX1 U60 ( .A(sfrwe), .Y(n44) );
  NOR32XL U61 ( .B(n227), .C(sfraddr[4]), .A(sfraddr[5]), .Y(n146) );
  NAND2X1 U62 ( .A(n181), .B(n87), .Y(n179) );
  NAND3X1 U63 ( .A(n193), .B(n17), .C(t_shift_clk), .Y(n176) );
  NAND4X1 U64 ( .A(sfraddr[0]), .B(sfraddr[4]), .C(n194), .D(n195), .Y(n193)
         );
  NOR4XL U65 ( .A(sfraddr[6]), .B(sfraddr[5]), .C(sfraddr[2]), .D(sfraddr[1]), 
        .Y(n195) );
  NOR2X1 U66 ( .A(n5), .B(n44), .Y(n194) );
  NAND41X1 U67 ( .D(sfraddr[4]), .A(sfraddr[5]), .B(n140), .C(n227), .Y(n228)
         );
  NAND4X1 U68 ( .A(sfraddr[5]), .B(n140), .C(sfraddr[4]), .D(n227), .Y(n226)
         );
  INVX1 U69 ( .A(sfraddr[3]), .Y(n5) );
  NOR3XL U70 ( .A(n25), .B(sfraddr[6]), .C(n4), .Y(n140) );
  INVX1 U71 ( .A(sfraddr[1]), .Y(n4) );
  INVX1 U72 ( .A(sfrdatai[5]), .Y(n11) );
  INVX1 U73 ( .A(sfrdatai[3]), .Y(n9) );
  INVX1 U74 ( .A(sfrdatai[4]), .Y(n10) );
  INVX1 U75 ( .A(sfrdatai[7]), .Y(n14) );
  INVX1 U76 ( .A(sfrdatai[2]), .Y(n8) );
  INVX1 U77 ( .A(sfrdatai[0]), .Y(n6) );
  INVX1 U78 ( .A(sfrdatai[6]), .Y(n12) );
  INVX1 U79 ( .A(sfrdatai[1]), .Y(n7) );
  NOR21XL U80 ( .B(t1ov), .A(n20), .Y(N59) );
  INVX1 U81 ( .A(n201), .Y(n47) );
  INVX1 U82 ( .A(n96), .Y(n45) );
  INVX1 U83 ( .A(n87), .Y(n51) );
  INVX1 U84 ( .A(rst), .Y(n30) );
  INVX1 U85 ( .A(rst), .Y(n31) );
  NAND2X1 U86 ( .A(n51), .B(n50), .Y(n112) );
  NAND2X1 U87 ( .A(n49), .B(n149), .Y(n147) );
  INVX1 U88 ( .A(rst), .Y(n29) );
  OAI222XL U89 ( .A(n40), .B(n6), .C(n113), .D(n252), .E(N108), .F(n253), .Y(
        n237) );
  OAI32X1 U90 ( .A(n73), .B(n23), .C(n34), .D(n139), .E(n14), .Y(n244) );
  INVX1 U91 ( .A(n139), .Y(n34) );
  NAND4X1 U92 ( .A(n140), .B(sfraddr[0]), .C(sfraddr[2]), .D(n141), .Y(n139)
         );
  NOR4XL U93 ( .A(sfraddr[5]), .B(sfraddr[4]), .C(sfraddr[3]), .D(n44), .Y(
        n141) );
  OAI32X1 U94 ( .A(n96), .B(n26), .C(n101), .D(n255), .E(n33), .Y(n232) );
  INVX1 U95 ( .A(n101), .Y(n33) );
  AOI221XL U96 ( .A(n96), .B(newinstr), .C(n97), .D(n45), .E(n28), .Y(n101) );
  GEN2XL U97 ( .D(n45), .E(n97), .C(n114), .B(n19), .A(n115), .Y(n238) );
  NOR4XL U98 ( .A(n23), .B(newinstr), .C(n45), .D(n252), .Y(n115) );
  NAND2X1 U99 ( .A(n52), .B(n53), .Y(n87) );
  NOR2X1 U100 ( .A(n87), .B(n74), .Y(rxd0oe) );
  AOI21BBXL U101 ( .B(n68), .C(n197), .A(n203), .Y(n201) );
  NAND4X1 U102 ( .A(r_shift_clk), .B(n98), .C(n87), .D(n253), .Y(n96) );
  NOR2X1 U103 ( .A(n128), .B(n22), .Y(n170) );
  INVX1 U104 ( .A(n128), .Y(n46) );
  OAI21X1 U105 ( .B(n71), .C(n121), .A(n18), .Y(n207) );
  AND3X1 U106 ( .A(n132), .B(n16), .C(n51), .Y(n162) );
  AOI22AXL U107 ( .A(n87), .B(n54), .D(n132), .C(n51), .Y(n150) );
  NAND4X1 U108 ( .A(n149), .B(r_shift_clk), .C(n112), .D(n253), .Y(n148) );
  AOI31X1 U109 ( .A(n161), .B(n154), .C(n3), .D(n162), .Y(n157) );
  NAND2X1 U110 ( .A(n98), .B(n100), .Y(n89) );
  OAI21X1 U111 ( .B(n27), .C(n130), .A(N382), .Y(n161) );
  INVX1 U112 ( .A(n221), .Y(n63) );
  OAI32X1 U113 ( .A(n70), .B(n121), .C(n207), .D(n208), .E(n71), .Y(N188) );
  OAI22X1 U114 ( .A(n147), .B(n86), .C(n148), .D(n246), .Y(N473) );
  OAI22X1 U115 ( .A(n147), .B(n85), .C(n148), .D(n86), .Y(N474) );
  OAI22X1 U116 ( .A(n147), .B(n84), .C(n148), .D(n85), .Y(N475) );
  OAI22X1 U117 ( .A(n147), .B(n83), .C(n148), .D(n84), .Y(N476) );
  OAI22X1 U118 ( .A(n147), .B(n82), .C(n148), .D(n83), .Y(N477) );
  OAI22X1 U119 ( .A(n81), .B(n147), .C(n148), .D(n82), .Y(N478) );
  OAI22X1 U120 ( .A(n76), .B(n147), .C(n148), .D(n81), .Y(N479) );
  NAND2X1 U121 ( .A(n128), .B(n15), .Y(N324) );
  OAI2B11X1 U122 ( .D(n97), .C(n148), .A(n147), .B(n17), .Y(N471) );
  NOR2X1 U123 ( .A(n74), .B(n131), .Y(t_shift_clk) );
  INVX1 U124 ( .A(n131), .Y(n50) );
  NAND2X1 U125 ( .A(n76), .B(n15), .Y(N382) );
  NOR2X1 U126 ( .A(n168), .B(n166), .Y(N363) );
  XNOR2XL U127 ( .A(n92), .B(n80), .Y(n168) );
  NAND3X1 U128 ( .A(n17), .B(n248), .C(n166), .Y(N360) );
  INVX1 U129 ( .A(n151), .Y(n13) );
  NAND2X1 U130 ( .A(n16), .B(n203), .Y(N223) );
  NAND2X1 U131 ( .A(n150), .B(n151), .Y(N428) );
  NOR21XL U132 ( .B(n98), .A(n21), .Y(n149) );
  NOR32XL U133 ( .B(n51), .C(n98), .A(n131), .Y(n114) );
  AOI21X1 U134 ( .B(n74), .C(n77), .A(n28), .Y(n116) );
  NAND32X1 U135 ( .B(n2), .C(n27), .A(n221), .Y(N166) );
  OAI21X1 U136 ( .B(n128), .C(n256), .A(n29), .Y(N325) );
  NOR2X1 U137 ( .A(n20), .B(n142), .Y(n245) );
  XNOR2XL U138 ( .A(n143), .B(n72), .Y(n142) );
  NAND2X1 U139 ( .A(n16), .B(n246), .Y(N375) );
  NAND2X1 U140 ( .A(n16), .B(n86), .Y(N376) );
  NAND2X1 U141 ( .A(n16), .B(n85), .Y(N377) );
  NAND2X1 U142 ( .A(n16), .B(n84), .Y(N378) );
  NAND2X1 U143 ( .A(n16), .B(n83), .Y(N379) );
  NAND2X1 U144 ( .A(n16), .B(n82), .Y(N380) );
  NAND2X1 U145 ( .A(n15), .B(n81), .Y(N381) );
  NOR3XL U146 ( .A(n222), .B(n25), .C(n206), .Y(N142) );
  NOR3XL U147 ( .A(n72), .B(n25), .C(n143), .Y(N207) );
  NOR2X1 U148 ( .A(n23), .B(n253), .Y(N348) );
  NOR2X1 U149 ( .A(n20), .B(n256), .Y(N307) );
  INVX1 U150 ( .A(n154), .Y(n54) );
  INVX1 U151 ( .A(n92), .Y(n79) );
  AO222X1 U152 ( .A(sfrdatai[1]), .B(n133), .C(ti_tmp), .D(n41), .E(s0con[1]), 
        .F(n39), .Y(n241) );
  OAI21X1 U153 ( .B(t_shift_count[0]), .C(n176), .A(n180), .Y(N281) );
  OAI21X1 U154 ( .B(s0con[7]), .C(n53), .A(n181), .Y(n180) );
  NAND3X1 U155 ( .A(n183), .B(n17), .C(n184), .Y(N267) );
  AOI22X1 U156 ( .A(t_shift_reg[10]), .B(n38), .C(sfrdatai[7]), .D(n181), .Y(
        n184) );
  OAI211X1 U157 ( .C(n6), .D(n179), .A(n18), .B(n191), .Y(N260) );
  AOI22X1 U158 ( .A(n36), .B(sfrdatai[1]), .C(t_shift_reg[3]), .D(n38), .Y(
        n191) );
  OAI211X1 U159 ( .C(n7), .D(n179), .A(n18), .B(n190), .Y(N261) );
  AOI22X1 U160 ( .A(n36), .B(sfrdatai[2]), .C(t_shift_reg[4]), .D(n38), .Y(
        n190) );
  OAI211X1 U161 ( .C(n179), .D(n11), .A(n18), .B(n186), .Y(N265) );
  AOI22X1 U162 ( .A(n36), .B(sfrdatai[6]), .C(t_shift_reg[8]), .D(n38), .Y(
        n186) );
  OAI211X1 U163 ( .C(n8), .D(n179), .A(n18), .B(n189), .Y(N262) );
  AOI22X1 U164 ( .A(sfrdatai[3]), .B(n36), .C(t_shift_reg[5]), .D(n38), .Y(
        n189) );
  OAI211X1 U165 ( .C(n40), .D(n8), .A(n93), .B(n94), .Y(n230) );
  NAND3X1 U166 ( .A(s0con2_tmp), .B(n41), .C(s0con2_val), .Y(n93) );
  NAND3X1 U167 ( .A(n39), .B(n255), .C(s0con[2]), .Y(n94) );
  OAI211X1 U168 ( .C(n179), .D(n9), .A(n18), .B(n188), .Y(N263) );
  AOI22X1 U169 ( .A(sfrdatai[4]), .B(n36), .C(t_shift_reg[6]), .D(n38), .Y(
        n188) );
  OAI211X1 U170 ( .C(n179), .D(n10), .A(n18), .B(n187), .Y(N264) );
  AOI22X1 U171 ( .A(sfrdatai[5]), .B(n36), .C(t_shift_reg[7]), .D(n38), .Y(
        n187) );
  OAI211X1 U172 ( .C(n179), .D(n12), .A(n18), .B(n185), .Y(N266) );
  AOI22X1 U173 ( .A(n36), .B(sfrdatai[7]), .C(t_shift_reg[9]), .D(n38), .Y(
        n185) );
  OAI211X1 U174 ( .C(n6), .D(n183), .A(n18), .B(n192), .Y(N259) );
  NAND2X1 U175 ( .A(t_shift_reg[2]), .B(n38), .Y(n192) );
  NAND3X1 U176 ( .A(n176), .B(n17), .C(n182), .Y(N268) );
  OAI21X1 U177 ( .B(s0con[3]), .C(n52), .A(n181), .Y(n182) );
  GEN2XL U178 ( .D(t_shift_count[1]), .E(t_shift_count[0]), .C(n178), .B(n38), 
        .A(n37), .Y(N282) );
  INVX1 U179 ( .A(n179), .Y(n37) );
  INVX1 U180 ( .A(n144), .Y(n42) );
  AOI32X1 U181 ( .A(bd), .B(n17), .C(n145), .D(sfrdatai[7]), .E(n43), .Y(n144)
         );
  INVX1 U182 ( .A(n145), .Y(n43) );
  NAND4XL U183 ( .A(sfraddr[6]), .B(n146), .C(n15), .D(n4), .Y(n145) );
  OAI21X1 U184 ( .B(n175), .C(n176), .A(n35), .Y(N284) );
  XOR2X1 U185 ( .A(n138), .B(t_shift_count[3]), .Y(n175) );
  OAI2B11X1 U186 ( .D(t_shift_reg[1]), .C(n176), .A(n35), .B(n17), .Y(N258) );
  AOI21X1 U187 ( .B(n138), .C(n177), .A(n176), .Y(N283) );
  NAND21X1 U188 ( .B(n178), .A(t_shift_count[2]), .Y(n177) );
  NAND2X1 U189 ( .A(n137), .B(n35), .Y(n243) );
  OAI211X1 U190 ( .C(t_shift_count[3]), .D(n138), .A(n18), .B(t_start), .Y(
        n137) );
  NOR2X1 U191 ( .A(n20), .B(n135), .Y(n242) );
  AOI32X1 U192 ( .A(t_shift_clk), .B(t_shift_count[0]), .C(n136), .D(ti_tmp), 
        .E(n32), .Y(n135) );
  NOR3XL U193 ( .A(t_shift_count[1]), .B(t_shift_count[3]), .C(
        t_shift_count[2]), .Y(n136) );
  INVX1 U194 ( .A(newinstr), .Y(n32) );
  INVX1 U195 ( .A(s0con[6]), .Y(n53) );
  INVX1 U196 ( .A(s0con[7]), .Y(n52) );
  INVX1 U197 ( .A(t_start), .Y(n74) );
  EORX1 U198 ( .A(baud_r2_clk), .B(n73), .C(n143), .D(n73), .Y(n128) );
  AOI21BBXL U199 ( .B(t_baud_count[1]), .C(n47), .A(N224), .Y(n199) );
  AND3X1 U200 ( .A(n100), .B(n46), .C(r_start), .Y(r_shift_clk) );
  NOR2X1 U201 ( .A(s0relh[7]), .B(r_clk_ov2), .Y(n206) );
  EORX1 U202 ( .A(t1ov_ff), .B(n204), .C(n204), .D(n205), .Y(n143) );
  NOR2X1 U203 ( .A(n53), .B(bd), .Y(n204) );
  AOI32X1 U204 ( .A(n65), .B(n53), .C(s0con[7]), .D(baud_rate_ov), .E(s0con[6]), .Y(n205) );
  INVX1 U205 ( .A(n206), .Y(n65) );
  NOR2X1 U206 ( .A(n47), .B(t_baud_count[0]), .Y(N224) );
  NAND2X1 U207 ( .A(n170), .B(t_start), .Y(n203) );
  ENOX1 U208 ( .A(n197), .B(n47), .C(n198), .D(t_baud_count[3]), .Y(N227) );
  OAI21X1 U209 ( .B(n47), .C(t_baud_count[2]), .A(n199), .Y(n198) );
  NOR21XL U210 ( .B(rxd0_fall_fl), .A(N324), .Y(n102) );
  AOI22X1 U211 ( .A(t_baud_ov), .B(n87), .C(clk_ov12), .D(n51), .Y(n131) );
  AOI21X1 U212 ( .B(n64), .C(r_clk_ov2), .A(n1), .Y(n211) );
  NOR41XL U213 ( .D(r_shift_count[0]), .A(r_shift_count[1]), .B(
        r_shift_count[2]), .C(r_shift_count[3]), .Y(n98) );
  AOI21BBXL U214 ( .B(clk_count[1]), .C(n207), .A(N185), .Y(n208) );
  GEN2XL U215 ( .D(n249), .E(n250), .C(n102), .B(fluctuation_conter[1]), .A(
        n103), .Y(n233) );
  INVX1 U216 ( .A(n104), .Y(n249) );
  NOR4XL U217 ( .A(fluctuation_conter[1]), .B(n102), .C(n104), .D(n250), .Y(
        n103) );
  OAI21X1 U218 ( .B(n90), .C(n68), .A(n163), .Y(n100) );
  NAND4X1 U219 ( .A(r_baud_count[3]), .B(n164), .C(n80), .D(n68), .Y(n163) );
  NAND2X1 U220 ( .A(rxd0_fall_fl), .B(n15), .Y(n104) );
  OAI33XL U221 ( .A(n254), .B(n26), .C(n95), .D(n76), .E(n28), .F(n96), .Y(
        n231) );
  INVX1 U222 ( .A(s0con2_val), .Y(n254) );
  NOR42XL U223 ( .C(n97), .D(n98), .A(n77), .B(n99), .Y(n95) );
  NAND3X1 U224 ( .A(n87), .B(n253), .C(n100), .Y(n99) );
  OAI32X1 U225 ( .A(n207), .B(clk_count[2]), .C(n121), .D(n208), .E(n70), .Y(
        N187) );
  OAI32X1 U226 ( .A(n104), .B(fluctuation_conter[0]), .C(n102), .D(n250), .E(
        n48), .Y(n234) );
  INVX1 U227 ( .A(n102), .Y(n48) );
  OAI32X1 U228 ( .A(n248), .B(n104), .C(n251), .D(n169), .E(n166), .Y(N362) );
  INVX1 U229 ( .A(fluctuation_conter[1]), .Y(n251) );
  AOI21X1 U230 ( .B(r_baud_count[1]), .C(n78), .A(n164), .Y(n169) );
  OAI32X1 U231 ( .A(n248), .B(n104), .C(n250), .D(r_baud_count[0]), .E(n166), 
        .Y(N361) );
  OAI32X1 U232 ( .A(n154), .B(n23), .C(n51), .D(n159), .E(n160), .Y(N425) );
  AOI21X1 U233 ( .B(r_shift_count[1]), .C(r_shift_count[0]), .A(n158), .Y(n159) );
  AOI21X1 U234 ( .B(n161), .C(n3), .A(n162), .Y(n160) );
  NAND41X1 U235 ( .D(n223), .A(tim_baud[8]), .B(tim_baud[9]), .C(n224), .Y(
        n222) );
  NAND3X1 U236 ( .A(tim_baud[6]), .B(tim_baud[5]), .C(tim_baud[7]), .Y(n223)
         );
  NOR32XL U237 ( .B(tim_baud[4]), .C(tim_baud[3]), .A(n225), .Y(n224) );
  NAND3X1 U238 ( .A(tim_baud[1]), .B(tim_baud[0]), .C(tim_baud[2]), .Y(n225)
         );
  NOR2X1 U239 ( .A(n78), .B(r_baud_count[1]), .Y(n164) );
  NAND3X1 U240 ( .A(r_start), .B(n248), .C(n170), .Y(n166) );
  NOR2X1 U241 ( .A(n207), .B(clk_count[0]), .Y(N185) );
  INVX1 U242 ( .A(r_baud_count[2]), .Y(n80) );
  OAI22AX1 U243 ( .D(r_shift_reg[0]), .C(n148), .A(n147), .B(n246), .Y(N472)
         );
  OAI21BX1 U244 ( .C(ri0_fall), .B(n109), .A(n110), .Y(n236) );
  NAND4X1 U245 ( .A(ri0_ff), .B(n109), .C(n15), .D(n253), .Y(n110) );
  OAI2B11X1 U246 ( .D(ri0_ff), .C(n111), .A(n112), .B(n17), .Y(n109) );
  NAND2X1 U247 ( .A(n51), .B(n253), .Y(n111) );
  OAI21X1 U248 ( .B(N382), .C(n152), .A(n153), .Y(N427) );
  GEN2XL U249 ( .D(n130), .E(n87), .C(n152), .B(n150), .A(n26), .Y(n153) );
  AOI21X1 U250 ( .B(n155), .C(r_shift_count[3]), .A(n108), .Y(n152) );
  OAI21X1 U251 ( .B(n199), .C(n75), .A(n200), .Y(N226) );
  NAND4X1 U252 ( .A(n201), .B(t_baud_count[1]), .C(t_baud_count[0]), .D(n75), 
        .Y(n200) );
  INVX1 U253 ( .A(t_baud_count[2]), .Y(n75) );
  OAI21X1 U254 ( .B(n77), .C(n123), .A(n124), .Y(n240) );
  OAI211X1 U255 ( .C(n108), .D(n125), .A(n123), .B(n19), .Y(n124) );
  NAND42X1 U256 ( .C(n125), .D(n114), .A(n126), .B(n15), .Y(n123) );
  NOR3XL U257 ( .A(n87), .B(r_start), .C(n132), .Y(n125) );
  INVX1 U258 ( .A(s0relh[6]), .Y(n68) );
  AOI21X1 U259 ( .B(n155), .C(n156), .A(n157), .Y(N426) );
  NAND21X1 U260 ( .B(n158), .A(r_shift_count[2]), .Y(n156) );
  NAND3X1 U261 ( .A(ri0_fall), .B(n50), .C(s0con[4]), .Y(n132) );
  NAND2X1 U262 ( .A(n127), .B(n3), .Y(n126) );
  ENOX1 U263 ( .A(n128), .B(n129), .C(n108), .D(n54), .Y(n127) );
  AOI31X1 U264 ( .A(rxd0_val), .B(n100), .C(n130), .D(n67), .Y(n129) );
  INVX1 U265 ( .A(n89), .Y(n67) );
  INVX1 U266 ( .A(r_baud_count[0]), .Y(n78) );
  NOR2X1 U267 ( .A(n165), .B(n166), .Y(N364) );
  XNOR2XL U268 ( .A(r_baud_count[3]), .B(n167), .Y(n165) );
  NOR2X1 U269 ( .A(n80), .B(n92), .Y(n167) );
  NOR2X1 U270 ( .A(n202), .B(n47), .Y(N225) );
  XNOR2XL U271 ( .A(t_baud_count[1]), .B(t_baud_count[0]), .Y(n202) );
  NOR2X1 U272 ( .A(r_shift_count[0]), .B(n157), .Y(N424) );
  NOR2X1 U273 ( .A(n23), .B(n217), .Y(N170) );
  AOI22X1 U274 ( .A(N148), .B(n211), .C(s0rell[3]), .D(n63), .Y(n217) );
  NOR2X1 U275 ( .A(n20), .B(n218), .Y(N169) );
  AOI22X1 U276 ( .A(N147), .B(n2), .C(s0rell[2]), .D(n63), .Y(n218) );
  NAND2X1 U277 ( .A(r_baud_count[2]), .B(n164), .Y(n90) );
  NOR4XL U278 ( .A(n196), .B(t_baud_count[1]), .C(t_baud_count[3]), .D(
        t_baud_count[2]), .Y(N230) );
  NAND2X1 U279 ( .A(t_baud_count[0]), .B(n170), .Y(n196) );
  INVX1 U280 ( .A(n212), .Y(n61) );
  AOI221XL U281 ( .A(s0relh[0]), .B(n63), .C(N153), .D(n211), .E(n27), .Y(n212) );
  INVX1 U282 ( .A(n213), .Y(n55) );
  AOI221XL U283 ( .A(s0rell[7]), .B(n63), .C(N152), .D(n211), .E(n26), .Y(n213) );
  INVX1 U284 ( .A(n214), .Y(n56) );
  AOI221XL U285 ( .A(s0rell[6]), .B(n63), .C(N151), .D(n211), .E(n27), .Y(n214) );
  INVX1 U286 ( .A(n215), .Y(n57) );
  AOI221XL U287 ( .A(s0rell[5]), .B(n63), .C(N150), .D(n211), .E(n26), .Y(n215) );
  INVX1 U288 ( .A(n216), .Y(n58) );
  AOI221XL U289 ( .A(s0rell[4]), .B(n63), .C(N149), .D(n211), .E(n27), .Y(n216) );
  INVX1 U290 ( .A(n219), .Y(n59) );
  AOI221XL U291 ( .A(s0rell[1]), .B(n63), .C(N146), .D(n211), .E(n26), .Y(n219) );
  INVX1 U292 ( .A(n220), .Y(n60) );
  AOI221XL U293 ( .A(s0rell[0]), .B(n63), .C(N145), .D(n211), .E(n26), .Y(n220) );
  INVX1 U294 ( .A(n210), .Y(n62) );
  AOI221XL U295 ( .A(s0relh[1]), .B(n63), .C(N154), .D(n211), .E(n27), .Y(n210) );
  AO44X1 U296 ( .A(rxd0_fall_fl), .B(n105), .C(n66), .D(n17), .E(n98), .F(
        s0con[6]), .G(rxd0_ff), .H(n106), .Y(n235) );
  INVX1 U297 ( .A(n107), .Y(n66) );
  NAND2X1 U298 ( .A(rxd0_fall), .B(n108), .Y(n105) );
  NOR4XL U299 ( .A(s0con[7]), .B(rxd0ff), .C(n27), .D(n107), .Y(n106) );
  NAND21X1 U300 ( .B(r_shift_count[2]), .A(n158), .Y(n155) );
  NOR42XL U301 ( .C(r_shift_count[3]), .D(r_shift_count[1]), .A(
        r_shift_count[0]), .B(r_shift_count[2]), .Y(n130) );
  AND2X1 U302 ( .A(clk_count[0]), .B(n16), .Y(N190) );
  OAI33XL U303 ( .A(n88), .B(n52), .C(n247), .D(n89), .E(n27), .F(n52), .Y(
        n229) );
  INVX1 U304 ( .A(receive_11_bits), .Y(n247) );
  OAI31XL U305 ( .A(n90), .B(s0relh[6]), .C(r_baud_count[3]), .D(n91), .Y(n88)
         );
  AOI31X1 U306 ( .A(s0relh[6]), .B(n80), .C(n79), .D(n24), .Y(n91) );
  NAND41X1 U307 ( .D(t_baud_count[3]), .A(t_baud_count[2]), .B(t_baud_count[1]), .C(t_baud_count[0]), .Y(n197) );
  NOR2X1 U308 ( .A(r_shift_count[1]), .B(r_shift_count[0]), .Y(n158) );
  NOR2X1 U309 ( .A(n155), .B(r_shift_count[3]), .Y(n108) );
  OAI21X1 U310 ( .B(n3), .C(n256), .A(n171), .Y(N333) );
  AOI21X1 U311 ( .B(n172), .C(n3), .A(n28), .Y(n171) );
  NOR42XL U312 ( .C(n70), .D(N190), .A(n71), .B(clk_count[1]), .Y(N191) );
  NOR2X1 U313 ( .A(n209), .B(n207), .Y(N186) );
  XNOR2XL U314 ( .A(clk_count[1]), .B(clk_count[0]), .Y(n209) );
  OAI21BBX1 U315 ( .A(n46), .B(rxd0_vec[1]), .C(n19), .Y(N327) );
  OAI21BBX1 U316 ( .A(n46), .B(rxd0_vec[0]), .C(n31), .Y(N326) );
  INVX1 U317 ( .A(smod), .Y(n73) );
  NAND3X1 U318 ( .A(n116), .B(n117), .C(n118), .Y(n239) );
  NAND4X1 U319 ( .A(t_shift_count[3]), .B(t_shift_count[0]), .C(txd0), .D(n122), .Y(n117) );
  AOI22X1 U320 ( .A(n51), .B(n119), .C(t_shift_reg[0]), .D(n3), .Y(n118) );
  NOR3XL U321 ( .A(n3), .B(t_shift_count[2]), .C(t_shift_count[1]), .Y(n122)
         );
  AOI22X1 U322 ( .A(n68), .B(r_baud_count[3]), .C(r_baud_count[2]), .D(
        s0relh[6]), .Y(n107) );
  NAND21X1 U323 ( .B(t_shift_count[2]), .A(n178), .Y(n138) );
  NAND32X1 U324 ( .B(t_shift_reg[0]), .C(n3), .A(n116), .Y(N303) );
  INVX1 U325 ( .A(s0con[0]), .Y(n253) );
  NAND2X1 U326 ( .A(r_baud_count[1]), .B(r_baud_count[0]), .Y(n92) );
  NAND2X1 U327 ( .A(clk_count[1]), .B(clk_count[0]), .Y(n121) );
  NAND2X1 U328 ( .A(s0con[4]), .B(rxd0_fall), .Y(n154) );
  NOR2X1 U329 ( .A(t_shift_count[1]), .B(t_shift_count[0]), .Y(n178) );
  INVX1 U330 ( .A(rxd0_val), .Y(n76) );
  OAI31XL U331 ( .A(n69), .B(clk_count[3]), .C(clk_count[2]), .D(n120), .Y(
        n119) );
  INVX1 U332 ( .A(n121), .Y(n69) );
  OAI31XL U333 ( .A(clk_count[0]), .B(clk_count[2]), .C(clk_count[1]), .D(
        clk_count[3]), .Y(n120) );
  NOR4XL U334 ( .A(n173), .B(receive_11_bits), .C(rxd0_fall), .D(n26), .Y(N306) );
  OAI21X1 U335 ( .B(n174), .C(rxd0_fall_fl), .A(n77), .Y(n173) );
  NOR21XL U337 ( .B(rxd0_ff), .A(rxd0ff), .Y(n174) );
  INVX1 U338 ( .A(r_start), .Y(n77) );
  NAND2X1 U339 ( .A(s0con[5]), .B(n76), .Y(n97) );
  INVX1 U340 ( .A(clk_count[3]), .Y(n71) );
  INVX1 U341 ( .A(s0relh[7]), .Y(n64) );
  INVX1 U342 ( .A(rxd0_fall), .Y(n248) );
  INVX1 U343 ( .A(rxd0ff), .Y(n256) );
  INVX1 U344 ( .A(fluctuation_conter[0]), .Y(n250) );
  INVX1 U345 ( .A(clk_count[2]), .Y(n70) );
  INVX1 U346 ( .A(r_shift_reg[7]), .Y(n81) );
  INVX1 U347 ( .A(r_shift_reg[1]), .Y(n246) );
  INVX1 U348 ( .A(r_shift_reg[2]), .Y(n86) );
  INVX1 U349 ( .A(r_shift_reg[3]), .Y(n85) );
  INVX1 U350 ( .A(r_shift_reg[4]), .Y(n84) );
  INVX1 U351 ( .A(r_shift_reg[5]), .Y(n83) );
  INVX1 U352 ( .A(r_shift_reg[6]), .Y(n82) );
  INVX1 U353 ( .A(ri_tmp), .Y(n252) );
  INVX1 U354 ( .A(baud_r_count), .Y(n72) );
  INVX1 U355 ( .A(s0con2_tmp), .Y(n255) );
endmodule


module serial0_a0_DW01_inc_0 ( A, SUM );
  input [9:0] A;
  output [9:0] SUM;

  wire   [9:2] carry;

  HAD1X1 U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .SO(SUM[8]) );
  HAD1X1 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .SO(SUM[7]) );
  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  XOR2X1 U1 ( .A(carry[9]), .B(A[9]), .Y(SUM[9]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_serial0_a0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_serial0_a0_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_serial0_a0_3 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_serial0_a0_4 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_serial0_a0_5 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_serial0_a0_6 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_serial0_a0_7 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_serial0_a0_8 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_serial0_a0_9 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_serial0_a0_10 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_serial0_a0_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module ports_a0 ( clkper, rst, port0, sfrdatai, sfraddr, sfrwe );
  output [7:0] port0;
  input [7:0] sfrdatai;
  input [6:0] sfraddr;
  input clkper, rst, sfrwe;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, net12328, n2, n3, n4, n1;

  SNPS_CLOCK_GATE_HIGH_ports_a0 clk_gate_p0_reg ( .CLK(clkper), .EN(N2), 
        .ENCLK(net12328), .TE(1'b0) );
  DFFQX1 p0_reg_2_ ( .D(N5), .C(net12328), .Q(port0[2]) );
  DFFQX1 p0_reg_7_ ( .D(N10), .C(net12328), .Q(port0[7]) );
  DFFQX1 p0_reg_6_ ( .D(N9), .C(net12328), .Q(port0[6]) );
  DFFQX1 p0_reg_5_ ( .D(N8), .C(net12328), .Q(port0[5]) );
  DFFQX1 p0_reg_4_ ( .D(N7), .C(net12328), .Q(port0[4]) );
  DFFQX1 p0_reg_1_ ( .D(N4), .C(net12328), .Q(port0[1]) );
  DFFQX1 p0_reg_3_ ( .D(N6), .C(net12328), .Q(port0[3]) );
  DFFQX1 p0_reg_0_ ( .D(N3), .C(net12328), .Q(port0[0]) );
  NAND2X1 U2 ( .A(n1), .B(n2), .Y(N2) );
  NAND42X1 U3 ( .C(sfraddr[3]), .D(sfraddr[2]), .A(n3), .B(n4), .Y(n2) );
  NOR3XL U4 ( .A(sfraddr[4]), .B(sfraddr[6]), .C(sfraddr[5]), .Y(n3) );
  NOR42XL U5 ( .C(sfrwe), .D(n1), .A(sfraddr[1]), .B(sfraddr[0]), .Y(n4) );
  NOR21XL U6 ( .B(sfrdatai[0]), .A(n2), .Y(N3) );
  NOR21XL U7 ( .B(sfrdatai[1]), .A(n2), .Y(N4) );
  NOR21XL U8 ( .B(sfrdatai[2]), .A(n2), .Y(N5) );
  NOR21XL U9 ( .B(sfrdatai[3]), .A(n2), .Y(N6) );
  NOR21XL U10 ( .B(sfrdatai[4]), .A(n2), .Y(N7) );
  NOR21XL U11 ( .B(sfrdatai[5]), .A(n2), .Y(N8) );
  NOR21XL U12 ( .B(sfrdatai[6]), .A(n2), .Y(N9) );
  NOR21XL U13 ( .B(sfrdatai[7]), .A(n2), .Y(N10) );
  INVX1 U14 ( .A(rst), .Y(n1) );
endmodule


module SNPS_CLOCK_GATE_HIGH_ports_a0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module mdu_a0 ( clkper, rst, mdubsy, sfrdatai, sfraddr, sfrwe, sfroe, arcon, 
        md0, md1, md2, md3, md4, md5 );
  input [7:0] sfrdatai;
  input [6:0] sfraddr;
  output [7:0] arcon;
  output [7:0] md0;
  output [7:0] md1;
  output [7:0] md2;
  output [7:0] md3;
  output [7:0] md4;
  output [7:0] md5;
  input clkper, rst, sfrwe, sfroe;
  output mdubsy;
  wire   N95, N96, N97, N98, N104, N105, N106, N107, N108, N109, setmdef, N190,
         N191, N192, N193, N194, N195, N196, N197, N198, N258, N259, N260,
         N261, N262, N263, N264, N265, N266, N332, N333, N334, N335, N336,
         N337, N338, N339, N340, N405, N406, N407, N408, N409, N410, N411,
         N412, N413, N453, N454, N455, N456, N457, N458, N459, N460, N461,
         N483, N484, N485, N486, N487, N488, N489, N490, N491, N566, N567,
         N568, N569, N570, N571, N572, N573, N574, N575, N576, N577, N578,
         N579, N580, N581, N610, N612, N613, N614, N674, N675, N676, N677,
         N678, set_div16, set_div32, N802, N892, N893, N894, N895, net12346,
         net12352, net12357, net12362, net12367, net12372, net12377, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
         n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
         n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238,
         n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249,
         n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
         n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271,
         n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
         n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n3,
         n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, SYNOPSYS_UNCONNECTED_1,
         SYNOPSYS_UNCONNECTED_2;
  wire   [3:0] oper_reg;
  wire   [4:1] counter_st;
  wire   [17:1] sum1;
  wire   [17:1] sum;
  wire   [15:0] norm_reg;
  wire   [1:0] mdu_op;
  wire   [17:0] arg_a;
  wire   [16:1] arg_b;
  wire   [17:0] arg_c;
  wire   [16:1] arg_d;
  wire   [4:3] r384_carry;

  SNPS_CLOCK_GATE_HIGH_mdu_a0_0 clk_gate_arcon_s_reg ( .CLK(clkper), .EN(N104), 
        .ENCLK(net12346), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mdu_a0_6 clk_gate_md0_s_reg ( .CLK(clkper), .EN(N190), 
        .ENCLK(net12352), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mdu_a0_5 clk_gate_md1_s_reg ( .CLK(clkper), .EN(N258), 
        .ENCLK(net12357), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mdu_a0_4 clk_gate_md2_s_reg ( .CLK(clkper), .EN(N332), 
        .ENCLK(net12362), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mdu_a0_3 clk_gate_md3_s_reg ( .CLK(clkper), .EN(N405), 
        .ENCLK(net12367), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mdu_a0_2 clk_gate_md4_s_reg ( .CLK(clkper), .EN(N453), 
        .ENCLK(net12372), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mdu_a0_1 clk_gate_md5_s_reg ( .CLK(clkper), .EN(N483), 
        .ENCLK(net12377), .TE(1'b0) );
  mdu_a0_DW01_add_0 add_1040 ( .A(arg_c), .B({1'b0, arg_d, n29}), .CI(1'b0), 
        .SUM({sum, SYNOPSYS_UNCONNECTED_1}), .CO() );
  mdu_a0_DW01_add_1 add_961 ( .A({arg_a[17:1], n30}), .B({1'b0, arg_b, n29}), 
        .CI(1'b0), .SUM({sum1, SYNOPSYS_UNCONNECTED_2}), .CO() );
  DFFQX1 setmdef_reg ( .D(N802), .C(clkper), .Q(setmdef) );
  DFFQX1 set_div16_reg ( .D(n414), .C(clkper), .Q(set_div16) );
  DFFQX1 set_div32_reg ( .D(n413), .C(clkper), .Q(set_div32) );
  DFFQX1 counter_st_reg_0_ ( .D(N674), .C(clkper), .Q(N610) );
  DFFQX1 counter_st_reg_2_ ( .D(N676), .C(clkper), .Q(counter_st[2]) );
  DFFQX1 counter_st_reg_4_ ( .D(N678), .C(clkper), .Q(counter_st[4]) );
  DFFQX1 counter_st_reg_3_ ( .D(N677), .C(clkper), .Q(counter_st[3]) );
  DFFQX1 counter_st_reg_1_ ( .D(N675), .C(clkper), .Q(counter_st[1]) );
  DFFQX1 oper_reg_reg_1_ ( .D(N893), .C(clkper), .Q(oper_reg[1]) );
  DFFQX1 oper_reg_reg_0_ ( .D(N892), .C(clkper), .Q(oper_reg[0]) );
  DFFQX1 oper_reg_reg_3_ ( .D(N895), .C(clkper), .Q(oper_reg[3]) );
  DFFQX1 oper_reg_reg_2_ ( .D(N894), .C(clkper), .Q(oper_reg[2]) );
  DFFQX1 norm_reg_reg_15_ ( .D(N581), .C(clkper), .Q(norm_reg[15]) );
  DFFQX1 norm_reg_reg_14_ ( .D(N580), .C(clkper), .Q(norm_reg[14]) );
  DFFQX1 norm_reg_reg_13_ ( .D(N579), .C(clkper), .Q(norm_reg[13]) );
  DFFQX1 norm_reg_reg_12_ ( .D(N578), .C(clkper), .Q(norm_reg[12]) );
  DFFQX1 norm_reg_reg_11_ ( .D(N577), .C(clkper), .Q(norm_reg[11]) );
  DFFQX1 norm_reg_reg_10_ ( .D(N576), .C(clkper), .Q(norm_reg[10]) );
  DFFQX1 norm_reg_reg_8_ ( .D(N574), .C(clkper), .Q(norm_reg[8]) );
  DFFQX1 norm_reg_reg_9_ ( .D(N575), .C(clkper), .Q(norm_reg[9]) );
  DFFQX1 arcon_s_reg_7_ ( .D(n410), .C(clkper), .Q(arcon[7]) );
  DFFQX1 arcon_s_reg_6_ ( .D(n408), .C(clkper), .Q(arcon[6]) );
  DFFQX1 arcon_s_reg_4_ ( .D(N109), .C(net12346), .Q(arcon[4]) );
  DFFQX1 md0_s_reg_2_ ( .D(N193), .C(net12352), .Q(md0[2]) );
  DFFQX1 norm_reg_reg_7_ ( .D(N573), .C(clkper), .Q(norm_reg[7]) );
  DFFQX1 arcon_s_reg_5_ ( .D(n409), .C(net12346), .Q(arcon[5]) );
  DFFQX1 md1_s_reg_5_ ( .D(N264), .C(net12357), .Q(md1[5]) );
  DFFQX1 md1_s_reg_6_ ( .D(N265), .C(net12357), .Q(md1[6]) );
  DFFQX1 md1_s_reg_4_ ( .D(N263), .C(net12357), .Q(md1[4]) );
  DFFQX1 md5_s_reg_7_ ( .D(N491), .C(net12377), .Q(md5[7]) );
  DFFQX1 md5_s_reg_6_ ( .D(N490), .C(net12377), .Q(md5[6]) );
  DFFQX1 md3_s_reg_2_ ( .D(N408), .C(net12367), .Q(md3[2]) );
  DFFQX1 md1_s_reg_2_ ( .D(N261), .C(net12357), .Q(md1[2]) );
  DFFQX1 md3_s_reg_6_ ( .D(N412), .C(net12367), .Q(md3[6]) );
  DFFQX1 md5_s_reg_2_ ( .D(N486), .C(net12377), .Q(md5[2]) );
  DFFQX1 arcon_s_reg_2_ ( .D(N107), .C(net12346), .Q(arcon[2]) );
  DFFQX1 arcon_s_reg_1_ ( .D(N106), .C(net12346), .Q(arcon[1]) );
  DFFQX1 arcon_s_reg_0_ ( .D(N105), .C(net12346), .Q(arcon[0]) );
  DFFQX1 arcon_s_reg_3_ ( .D(N108), .C(net12346), .Q(arcon[3]) );
  DFFQX1 md0_s_reg_1_ ( .D(N192), .C(net12352), .Q(md0[1]) );
  DFFQX1 norm_reg_reg_6_ ( .D(N572), .C(clkper), .Q(norm_reg[6]) );
  DFFQX1 norm_reg_reg_5_ ( .D(N571), .C(clkper), .Q(norm_reg[5]) );
  DFFQX1 md1_s_reg_0_ ( .D(N259), .C(net12357), .Q(md1[0]) );
  DFFQX1 md3_s_reg_4_ ( .D(N410), .C(net12367), .Q(md3[4]) );
  DFFQX1 md0_s_reg_3_ ( .D(N194), .C(net12352), .Q(md0[3]) );
  DFFQX1 md1_s_reg_1_ ( .D(N260), .C(net12357), .Q(md1[1]) );
  DFFQX1 md1_s_reg_3_ ( .D(N262), .C(net12357), .Q(md1[3]) );
  DFFQX1 md0_s_reg_4_ ( .D(N195), .C(net12352), .Q(md0[4]) );
  DFFQX1 md0_s_reg_5_ ( .D(N196), .C(net12352), .Q(md0[5]) );
  DFFQX1 md0_s_reg_6_ ( .D(N197), .C(net12352), .Q(md0[6]) );
  DFFQX1 md0_s_reg_7_ ( .D(N198), .C(net12352), .Q(md0[7]) );
  DFFQX1 md5_s_reg_3_ ( .D(N487), .C(net12377), .Q(md5[3]) );
  DFFQX1 md4_s_reg_6_ ( .D(N460), .C(net12372), .Q(md4[6]) );
  DFFQX1 md5_s_reg_4_ ( .D(N488), .C(net12377), .Q(md5[4]) );
  DFFQX1 md3_s_reg_1_ ( .D(N407), .C(net12367), .Q(md3[1]) );
  DFFQX1 md3_s_reg_0_ ( .D(N406), .C(net12367), .Q(md3[0]) );
  DFFQX1 md2_s_reg_7_ ( .D(N340), .C(net12362), .Q(md2[7]) );
  DFFQX1 md5_s_reg_5_ ( .D(N489), .C(net12377), .Q(md5[5]) );
  DFFQX1 md3_s_reg_3_ ( .D(N409), .C(net12367), .Q(md3[3]) );
  DFFQX1 md5_s_reg_1_ ( .D(N485), .C(net12377), .Q(md5[1]) );
  DFFQX1 md4_s_reg_7_ ( .D(N461), .C(net12372), .Q(md4[7]) );
  DFFQX1 md3_s_reg_5_ ( .D(N411), .C(net12367), .Q(md3[5]) );
  DFFQX1 md5_s_reg_0_ ( .D(N484), .C(net12377), .Q(md5[0]) );
  DFFQX1 norm_reg_reg_4_ ( .D(N570), .C(clkper), .Q(norm_reg[4]) );
  DFFQX1 md4_s_reg_5_ ( .D(N459), .C(net12372), .Q(md4[5]) );
  DFFQX1 md2_s_reg_5_ ( .D(N338), .C(net12362), .Q(md2[5]) );
  DFFQX1 md2_s_reg_6_ ( .D(N339), .C(net12362), .Q(md2[6]) );
  DFFQX1 norm_reg_reg_2_ ( .D(N568), .C(clkper), .Q(norm_reg[2]) );
  DFFQX1 norm_reg_reg_3_ ( .D(N569), .C(clkper), .Q(norm_reg[3]) );
  DFFQX1 md4_s_reg_4_ ( .D(N458), .C(net12372), .Q(md4[4]) );
  DFFQX1 md4_s_reg_3_ ( .D(N457), .C(net12372), .Q(md4[3]) );
  DFFQX1 md2_s_reg_4_ ( .D(N337), .C(net12362), .Q(md2[4]) );
  DFFQX1 md2_s_reg_3_ ( .D(N336), .C(net12362), .Q(md2[3]) );
  DFFQX1 norm_reg_reg_1_ ( .D(N567), .C(clkper), .Q(norm_reg[1]) );
  DFFQX1 md4_s_reg_2_ ( .D(N456), .C(net12372), .Q(md4[2]) );
  DFFQX1 md2_s_reg_2_ ( .D(N335), .C(net12362), .Q(md2[2]) );
  DFFQX1 norm_reg_reg_0_ ( .D(N566), .C(clkper), .Q(norm_reg[0]) );
  DFFQX1 md2_s_reg_0_ ( .D(N333), .C(net12362), .Q(md2[0]) );
  DFFQX1 md2_s_reg_1_ ( .D(N334), .C(net12362), .Q(md2[1]) );
  DFFQX1 md4_s_reg_0_ ( .D(N454), .C(net12372), .Q(md4[0]) );
  DFFQX1 md4_s_reg_1_ ( .D(N455), .C(net12372), .Q(md4[1]) );
  DFFQX1 md0_s_reg_0_ ( .D(N191), .C(net12352), .Q(md0[0]) );
  DFFQX1 md1_s_reg_7_ ( .D(N266), .C(net12357), .Q(md1[7]) );
  DFFQX1 md3_s_reg_7_ ( .D(N413), .C(net12367), .Q(md3[7]) );
  DFFQX1 mdu_op_reg_0_ ( .D(n411), .C(clkper), .Q(mdu_op[0]) );
  DFFQX1 mdu_op_reg_1_ ( .D(n412), .C(clkper), .Q(mdu_op[1]) );
  INVX1 U3 ( .A(n53), .Y(n3) );
  INVX1 U4 ( .A(n384), .Y(n4) );
  NAND2X1 U5 ( .A(n277), .B(n74), .Y(n5) );
  INVX1 U6 ( .A(n303), .Y(n6) );
  NAND2X1 U7 ( .A(arg_c[0]), .B(n68), .Y(n7) );
  BUFX3 U8 ( .A(n258), .Y(n8) );
  NAND2X1 U9 ( .A(n18), .B(n108), .Y(n9) );
  INVX1 U10 ( .A(n106), .Y(n10) );
  INVX1 U11 ( .A(n300), .Y(n11) );
  NAND2X1 U12 ( .A(sum1[17]), .B(arg_c[0]), .Y(n12) );
  BUFX3 U13 ( .A(n199), .Y(n13) );
  BUFX3 U14 ( .A(n262), .Y(n14) );
  BUFX3 U15 ( .A(n347), .Y(n15) );
  INVX1 U16 ( .A(n302), .Y(n16) );
  BUFX3 U17 ( .A(n193), .Y(n17) );
  NOR2X1 U18 ( .A(sum1[17]), .B(sum[17]), .Y(n18) );
  INVX1 U19 ( .A(n179), .Y(n19) );
  BUFX3 U20 ( .A(n306), .Y(n20) );
  INVX1 U21 ( .A(sum[17]), .Y(n23) );
  INVX1 U22 ( .A(n23), .Y(n21) );
  INVX1 U23 ( .A(n23), .Y(n22) );
  NOR4XL U24 ( .A(counter_st[1]), .B(counter_st[2]), .C(counter_st[3]), .D(
        counter_st[4]), .Y(n336) );
  NOR3XL U25 ( .A(n73), .B(n77), .C(n76), .Y(n245) );
  INVX1 U28 ( .A(n317), .Y(n73) );
  INVX1 U29 ( .A(n364), .Y(n76) );
  INVX1 U30 ( .A(n339), .Y(n77) );
  NOR2X1 U31 ( .A(n75), .B(n74), .Y(n242) );
  INVX1 U32 ( .A(n386), .Y(n75) );
  AOI21X1 U33 ( .B(n109), .C(n267), .A(n291), .Y(n338) );
  INVX1 U34 ( .A(n299), .Y(n24) );
  INVX1 U35 ( .A(n299), .Y(n25) );
  INVX1 U36 ( .A(n337), .Y(n105) );
  INVX1 U37 ( .A(n384), .Y(n100) );
  INVX1 U38 ( .A(n382), .Y(n103) );
  NOR32XL U39 ( .B(n338), .C(n340), .A(n341), .Y(n318) );
  AND3X1 U40 ( .A(n388), .B(n296), .C(n337), .Y(n340) );
  INVX1 U41 ( .A(n264), .Y(n108) );
  INVX1 U42 ( .A(n291), .Y(n98) );
  AOI21X1 U43 ( .B(n48), .C(n364), .A(n233), .Y(n190) );
  AOI21X1 U44 ( .B(n47), .C(n231), .A(n233), .Y(n268) );
  AOI21X1 U45 ( .B(n47), .C(n317), .A(n233), .Y(n292) );
  AOI21X1 U46 ( .B(n47), .C(n339), .A(n233), .Y(n319) );
  AOI21X1 U47 ( .B(n48), .C(n386), .A(n233), .Y(n368) );
  NAND2X1 U48 ( .A(n277), .B(n74), .Y(n185) );
  AOI31X1 U49 ( .A(n231), .B(n47), .C(n232), .D(n233), .Y(n201) );
  OAI21X1 U50 ( .B(n242), .C(n70), .A(n243), .Y(n189) );
  NAND2X1 U51 ( .A(n241), .B(n46), .Y(n191) );
  NAND2X1 U52 ( .A(n73), .B(n277), .Y(n186) );
  NAND2X1 U53 ( .A(n77), .B(n277), .Y(n187) );
  NAND2X1 U54 ( .A(n76), .B(n277), .Y(n345) );
  NAND2X1 U55 ( .A(n75), .B(n277), .Y(n367) );
  INVX1 U56 ( .A(n179), .Y(n71) );
  NOR2X1 U57 ( .A(n246), .B(n70), .Y(n241) );
  NAND3X1 U58 ( .A(n243), .B(n46), .C(n255), .Y(n391) );
  INVX1 U59 ( .A(n285), .Y(n69) );
  NAND4X1 U60 ( .A(n391), .B(n390), .C(n71), .D(n46), .Y(N104) );
  NAND2X1 U61 ( .A(n185), .B(n46), .Y(n183) );
  NAND3X1 U62 ( .A(n191), .B(n46), .C(n98), .Y(N453) );
  NAND3X1 U63 ( .A(n5), .B(n46), .C(n98), .Y(N483) );
  NAND3X1 U64 ( .A(n187), .B(n47), .C(n318), .Y(N332) );
  NAND3X1 U65 ( .A(n186), .B(n47), .C(n318), .Y(N405) );
  NAND3X1 U66 ( .A(n367), .B(n47), .C(n365), .Y(N190) );
  NAND3X1 U67 ( .A(n345), .B(n47), .C(n365), .Y(N258) );
  AND2X1 U68 ( .A(n366), .B(sfraddr[2]), .Y(n278) );
  NAND2X1 U69 ( .A(n344), .B(sfraddr[0]), .Y(n339) );
  NAND2X1 U70 ( .A(n344), .B(n35), .Y(n364) );
  NAND3X1 U71 ( .A(n35), .B(n36), .C(n278), .Y(n317) );
  INVX1 U72 ( .A(sfraddr[2]), .Y(n37) );
  NAND4X1 U73 ( .A(sfraddr[0]), .B(n366), .C(n36), .D(n37), .Y(n386) );
  INVX1 U74 ( .A(sfraddr[0]), .Y(n35) );
  NAND3X1 U75 ( .A(n278), .B(n36), .C(sfraddr[0]), .Y(n246) );
  INVX1 U76 ( .A(n232), .Y(n72) );
  INVX1 U77 ( .A(n231), .Y(n74) );
  NOR3XL U78 ( .A(n107), .B(n109), .C(n342), .Y(n291) );
  INVX1 U79 ( .A(n343), .Y(n107) );
  NAND2X1 U80 ( .A(n387), .B(n342), .Y(n388) );
  NAND3X1 U81 ( .A(n107), .B(n342), .C(n109), .Y(n337) );
  NOR2X1 U82 ( .A(n263), .B(n107), .Y(n387) );
  NAND3X1 U83 ( .A(n342), .B(n263), .C(n343), .Y(n296) );
  INVX1 U84 ( .A(n263), .Y(n109) );
  INVX1 U85 ( .A(n299), .Y(n101) );
  NOR21XL U86 ( .B(n387), .A(n342), .Y(n341) );
  NAND21X1 U87 ( .B(n341), .A(n306), .Y(n384) );
  NOR2X1 U88 ( .A(n342), .B(n387), .Y(n382) );
  NOR2X1 U89 ( .A(n342), .B(n343), .Y(n267) );
  NAND2X1 U90 ( .A(n342), .B(n263), .Y(n396) );
  INVX1 U91 ( .A(n255), .Y(n112) );
  NAND2X1 U92 ( .A(n267), .B(n46), .Y(n264) );
  NAND2X1 U93 ( .A(n262), .B(n108), .Y(n256) );
  NAND2X1 U94 ( .A(n18), .B(n108), .Y(n257) );
  NOR2X1 U95 ( .A(n14), .B(n259), .Y(n265) );
  INVX1 U96 ( .A(n34), .Y(n30) );
  INVX1 U97 ( .A(n29), .Y(n28) );
  INVX1 U98 ( .A(n33), .Y(n32) );
  NAND2X1 U99 ( .A(arg_c[0]), .B(n68), .Y(n195) );
  INVX1 U100 ( .A(n29), .Y(n26) );
  INVX1 U101 ( .A(n33), .Y(n31) );
  INVX1 U102 ( .A(n29), .Y(n27) );
  INVX1 U103 ( .A(sfrwe), .Y(n70) );
  NAND31X1 U104 ( .C(n406), .A(n46), .B(n243), .Y(n390) );
  NOR2X1 U105 ( .A(n241), .B(rst), .Y(n285) );
  NOR2X1 U106 ( .A(n70), .B(rst), .Y(n277) );
  NOR2X1 U107 ( .A(n243), .B(rst), .Y(n179) );
  NOR2XL U108 ( .A(rst), .B(sfrwe), .Y(n233) );
  NAND2XL U109 ( .A(sfrwe), .B(n72), .Y(n243) );
  AOI211X1 U110 ( .C(n238), .D(n239), .A(n240), .B(rst), .Y(N802) );
  EORX1 U111 ( .A(sfroe), .B(n244), .C(n245), .D(n70), .Y(n238) );
  NOR2X1 U112 ( .A(n241), .B(n189), .Y(n239) );
  NAND3X1 U113 ( .A(n245), .B(n246), .C(n242), .Y(n244) );
  AND3X1 U114 ( .A(n366), .B(n37), .C(sfraddr[1]), .Y(n344) );
  NOR43XL U115 ( .B(sfraddr[5]), .C(sfraddr[3]), .D(sfraddr[6]), .A(sfraddr[4]), .Y(n366) );
  NAND3X1 U116 ( .A(n278), .B(n35), .C(sfraddr[1]), .Y(n231) );
  NAND3X1 U117 ( .A(sfraddr[0]), .B(n278), .C(sfraddr[1]), .Y(n232) );
  INVX1 U118 ( .A(sfraddr[1]), .Y(n36) );
  INVX1 U119 ( .A(sfrdatai[4]), .Y(n42) );
  INVX1 U120 ( .A(sfrdatai[5]), .Y(n43) );
  INVX1 U121 ( .A(sfrdatai[3]), .Y(n41) );
  INVX1 U122 ( .A(sfrdatai[2]), .Y(n40) );
  INVX1 U123 ( .A(sfrdatai[1]), .Y(n39) );
  INVX1 U124 ( .A(sfrdatai[0]), .Y(n38) );
  INVX1 U125 ( .A(sfrdatai[7]), .Y(n45) );
  INVX1 U126 ( .A(sfrdatai[6]), .Y(n44) );
  NOR32XL U127 ( .B(n401), .C(n227), .A(n254), .Y(n343) );
  NAND4X1 U128 ( .A(n401), .B(n112), .C(n206), .D(n167), .Y(n342) );
  NAND2X1 U129 ( .A(n398), .B(n206), .Y(n263) );
  NOR2X1 U130 ( .A(n421), .B(n388), .Y(n299) );
  NOR42XL U131 ( .C(n401), .D(n212), .A(n110), .B(n166), .Y(n398) );
  INVX1 U132 ( .A(n300), .Y(n104) );
  INVX1 U133 ( .A(n351), .Y(n106) );
  INVX1 U134 ( .A(n167), .Y(n110) );
  INVX1 U135 ( .A(n302), .Y(n102) );
  NAND2X1 U136 ( .A(n235), .B(n227), .Y(n255) );
  NAND3X1 U137 ( .A(n212), .B(n206), .C(n210), .Y(n254) );
  NAND21X1 U138 ( .B(n388), .A(n421), .Y(n306) );
  AND4X1 U139 ( .A(n398), .B(n112), .C(n210), .D(n214), .Y(n394) );
  AND3X1 U140 ( .A(n302), .B(n340), .C(n103), .Y(n365) );
  OAI31XL U141 ( .A(n253), .B(n254), .C(n255), .D(n47), .Y(n248) );
  NAND2X1 U142 ( .A(n214), .B(n167), .Y(n253) );
  INVX1 U143 ( .A(rst), .Y(n46) );
  INVX1 U144 ( .A(rst), .Y(n47) );
  OAI22X1 U145 ( .A(n209), .B(n210), .C(n218), .D(n227), .Y(n225) );
  INVX1 U146 ( .A(rst), .Y(n48) );
  INVX1 U147 ( .A(n206), .Y(n113) );
  INVX1 U148 ( .A(n214), .Y(n115) );
  NOR2X1 U149 ( .A(sum1[17]), .B(sum[17]), .Y(n259) );
  NOR2X1 U150 ( .A(n68), .B(n22), .Y(n262) );
  NAND2X1 U151 ( .A(sum1[17]), .B(arg_c[0]), .Y(n194) );
  OAI222XL U152 ( .A(n80), .B(n256), .C(n431), .D(n257), .E(n258), .F(n54), 
        .Y(N581) );
  OAI222XL U153 ( .A(n82), .B(n256), .C(n430), .D(n9), .E(n258), .F(n56), .Y(
        N579) );
  INVX1 U154 ( .A(sum[14]), .Y(n56) );
  OAI222XL U155 ( .A(n84), .B(n256), .C(n429), .D(n257), .E(n258), .F(n58), 
        .Y(N577) );
  INVX1 U156 ( .A(sum[12]), .Y(n58) );
  OAI222XL U157 ( .A(n86), .B(n256), .C(n428), .D(n9), .E(n258), .F(n60), .Y(
        N575) );
  INVX1 U158 ( .A(sum[10]), .Y(n60) );
  OAI222XL U159 ( .A(n88), .B(n256), .C(n427), .D(n257), .E(n258), .F(n62), 
        .Y(N573) );
  INVX1 U160 ( .A(sum[8]), .Y(n62) );
  OAI222XL U161 ( .A(n90), .B(n256), .C(n426), .D(n9), .E(n258), .F(n64), .Y(
        N571) );
  INVX1 U162 ( .A(sum[6]), .Y(n64) );
  OAI222XL U163 ( .A(n92), .B(n256), .C(n425), .D(n257), .E(n258), .F(n66), 
        .Y(N569) );
  INVX1 U164 ( .A(sum[4]), .Y(n66) );
  OAI222XL U165 ( .A(n81), .B(n256), .C(n159), .D(n9), .E(n258), .F(n55), .Y(
        N580) );
  INVX1 U166 ( .A(sum[15]), .Y(n55) );
  OAI222XL U167 ( .A(n83), .B(n256), .C(n158), .D(n257), .E(n258), .F(n57), 
        .Y(N578) );
  INVX1 U168 ( .A(sum[13]), .Y(n57) );
  OAI222XL U169 ( .A(n85), .B(n3), .C(n157), .D(n9), .E(n8), .F(n59), .Y(N576)
         );
  INVX1 U170 ( .A(sum[11]), .Y(n59) );
  OAI222XL U171 ( .A(n87), .B(n3), .C(n156), .D(n257), .E(n8), .F(n61), .Y(
        N574) );
  INVX1 U172 ( .A(sum[9]), .Y(n61) );
  OAI222XL U173 ( .A(n89), .B(n3), .C(n155), .D(n9), .E(n8), .F(n63), .Y(N572)
         );
  INVX1 U174 ( .A(sum[7]), .Y(n63) );
  OAI222XL U175 ( .A(n91), .B(n3), .C(n154), .D(n257), .E(n8), .F(n65), .Y(
        N570) );
  INVX1 U176 ( .A(sum[5]), .Y(n65) );
  OAI222XL U177 ( .A(n94), .B(n3), .C(n146), .D(n9), .E(n8), .F(n67), .Y(N568)
         );
  INVX1 U178 ( .A(sum[3]), .Y(n67) );
  OAI21X1 U179 ( .B(n191), .C(n38), .A(n289), .Y(N454) );
  AOI33X1 U180 ( .A(n290), .B(n52), .C(n285), .D(sum[1]), .E(n21), .F(n285), 
        .Y(n289) );
  OAI22X1 U181 ( .A(n200), .B(n138), .C(n96), .D(n137), .Y(n290) );
  INVX1 U182 ( .A(n265), .Y(n52) );
  OAI21BX1 U183 ( .C(sum[2]), .B(n8), .A(n260), .Y(N567) );
  AOI32X1 U184 ( .A(n108), .B(n261), .C(n259), .D(n53), .E(sum1[1]), .Y(n260)
         );
  OAI22X1 U185 ( .A(n109), .B(n129), .C(n148), .D(n263), .Y(n261) );
  INVX1 U186 ( .A(n256), .Y(n53) );
  OAI21X1 U187 ( .B(n191), .C(n39), .A(n286), .Y(N455) );
  AOI32X1 U188 ( .A(n18), .B(n287), .C(n285), .D(n285), .E(n288), .Y(n286) );
  OAI22X1 U189 ( .A(n200), .B(n129), .C(n96), .D(n148), .Y(n287) );
  AO22X1 U190 ( .A(sum1[1]), .B(n14), .C(n21), .D(sum[2]), .Y(n288) );
  INVX1 U191 ( .A(n192), .Y(n29) );
  INVX1 U192 ( .A(arg_a[0]), .Y(n33) );
  INVX1 U193 ( .A(arg_a[0]), .Y(n34) );
  INVX1 U194 ( .A(sum[16]), .Y(n54) );
  NAND2X1 U195 ( .A(n22), .B(n108), .Y(n258) );
  INVX1 U196 ( .A(sum1[17]), .Y(n68) );
  OAI222XL U197 ( .A(N95), .B(n390), .C(n251), .D(n391), .E(n19), .F(n39), .Y(
        N106) );
  OAI222XL U198 ( .A(N96), .B(n390), .C(n250), .D(n391), .E(n71), .F(n40), .Y(
        N107) );
  OAI222XL U199 ( .A(N98), .B(n390), .C(n247), .D(n391), .E(n71), .F(n42), .Y(
        N109) );
  OAI222XL U200 ( .A(N97), .B(n390), .C(n249), .D(n391), .E(n71), .F(n41), .Y(
        N108) );
  OAI222XL U201 ( .A(n150), .B(n390), .C(n252), .D(n391), .E(n71), .F(n38), 
        .Y(N105) );
  OAI32X1 U202 ( .A(n116), .B(rst), .C(n179), .D(n71), .E(n43), .Y(n409) );
  OAI221X1 U203 ( .A(n185), .B(n78), .C(n183), .D(n97), .E(n71), .Y(n412) );
  OAI211X1 U204 ( .C(n201), .D(n202), .A(n185), .B(n71), .Y(N895) );
  AOI211X1 U205 ( .C(n110), .D(n203), .A(n204), .B(n205), .Y(n202) );
  OAI32X1 U206 ( .A(n206), .B(n148), .C(n207), .D(n29), .E(n208), .Y(n205) );
  OAI222XL U207 ( .A(n209), .B(n210), .C(n211), .D(n212), .E(n213), .F(n214), 
        .Y(n204) );
  AOI31X1 U208 ( .A(n229), .B(n111), .C(n230), .D(n201), .Y(N892) );
  INVX1 U209 ( .A(n226), .Y(n111) );
  OA22X1 U210 ( .A(n235), .B(n218), .C(n214), .D(n213), .Y(n229) );
  OA222X1 U211 ( .A(n212), .B(n151), .C(n219), .D(n116), .E(n208), .F(n200), 
        .Y(n230) );
  INVX1 U212 ( .A(sum1[2]), .Y(n94) );
  INVX1 U213 ( .A(sum1[4]), .Y(n91) );
  INVX1 U214 ( .A(sum1[5]), .Y(n90) );
  INVX1 U215 ( .A(sum1[6]), .Y(n89) );
  INVX1 U216 ( .A(sum1[7]), .Y(n88) );
  INVX1 U217 ( .A(sum1[8]), .Y(n87) );
  INVX1 U218 ( .A(sum1[9]), .Y(n86) );
  INVX1 U219 ( .A(sum1[10]), .Y(n85) );
  INVX1 U220 ( .A(sum1[11]), .Y(n84) );
  INVX1 U221 ( .A(sum1[12]), .Y(n83) );
  INVX1 U222 ( .A(sum1[13]), .Y(n82) );
  INVX1 U223 ( .A(sum1[14]), .Y(n81) );
  INVX1 U224 ( .A(sum1[15]), .Y(n80) );
  INVX1 U225 ( .A(sum1[3]), .Y(n92) );
  NAND2X1 U226 ( .A(n197), .B(n96), .Y(arg_c[0]) );
  INVX1 U227 ( .A(n200), .Y(n96) );
  OAI22X1 U228 ( .A(n421), .B(n337), .C(n137), .D(n296), .Y(n351) );
  NOR43XL U229 ( .B(n208), .C(n406), .D(n407), .A(n240), .Y(n401) );
  NOR21XL U230 ( .B(n171), .A(n161), .Y(n407) );
  OAI21X1 U231 ( .B(n137), .C(n296), .A(n297), .Y(n300) );
  NAND2X1 U232 ( .A(n403), .B(n404), .Y(n167) );
  OAI21X1 U233 ( .B(n336), .C(n337), .A(n338), .Y(n294) );
  AND2X1 U234 ( .A(n389), .B(n402), .Y(n161) );
  OAI31XL U235 ( .A(n149), .B(n152), .C(n117), .D(mdubsy), .Y(n240) );
  NAND2X1 U236 ( .A(n399), .B(n405), .Y(mdubsy) );
  NOR2X1 U237 ( .A(n114), .B(n117), .Y(n404) );
  NAND2X1 U238 ( .A(n399), .B(n404), .Y(n212) );
  NOR21XL U239 ( .B(n395), .A(n394), .Y(n393) );
  OAI211X1 U240 ( .C(n396), .D(n137), .A(n297), .B(n24), .Y(n395) );
  NAND2X1 U241 ( .A(n105), .B(n336), .Y(n297) );
  NOR2X1 U242 ( .A(n249), .B(n248), .Y(N677) );
  NOR2X1 U243 ( .A(n247), .B(n248), .Y(N678) );
  NOR2X1 U244 ( .A(n250), .B(n248), .Y(N676) );
  NOR2X1 U245 ( .A(n251), .B(n248), .Y(N675) );
  NOR2X1 U246 ( .A(n252), .B(n248), .Y(N674) );
  NAND2X1 U247 ( .A(n404), .B(n402), .Y(n406) );
  NAND2X1 U248 ( .A(n402), .B(n405), .Y(n171) );
  NAND2X1 U249 ( .A(n399), .B(n389), .Y(n206) );
  INVX1 U250 ( .A(n303), .Y(n99) );
  AND2X1 U251 ( .A(n400), .B(n402), .Y(n166) );
  AOI31X1 U252 ( .A(n397), .B(n20), .C(n342), .D(n394), .Y(n392) );
  AOI22AXL U253 ( .A(n421), .B(n105), .D(n396), .C(n137), .Y(n397) );
  NAND2X1 U254 ( .A(n341), .B(n223), .Y(n302) );
  NAND2X1 U255 ( .A(n403), .B(n405), .Y(n210) );
  NAND2X1 U256 ( .A(n403), .B(n400), .Y(n227) );
  NAND2X1 U257 ( .A(n403), .B(n389), .Y(n235) );
  INVX1 U258 ( .A(n336), .Y(n421) );
  NAND2X1 U259 ( .A(n399), .B(n400), .Y(n214) );
  GEN2XL U260 ( .D(n161), .E(n162), .C(n163), .B(n48), .A(n164), .Y(n408) );
  NAND4X1 U261 ( .A(n174), .B(n175), .C(n176), .D(n177), .Y(n162) );
  NOR4XL U262 ( .A(n165), .B(n166), .C(rst), .D(n161), .Y(n164) );
  OAI31XL U263 ( .A(n168), .B(n169), .C(n170), .D(n171), .Y(n163) );
  NAND2X1 U264 ( .A(n228), .B(n423), .Y(n209) );
  NAND2X1 U265 ( .A(n113), .B(n207), .Y(n219) );
  NAND2X1 U266 ( .A(n421), .B(n237), .Y(n218) );
  NAND4X1 U267 ( .A(n150), .B(n422), .C(n424), .D(n423), .Y(n237) );
  NAND4X1 U268 ( .A(n166), .B(n153), .C(n439), .D(n147), .Y(n170) );
  INVX1 U269 ( .A(n211), .Y(n151) );
  AND3X1 U270 ( .A(n178), .B(n130), .C(n139), .Y(n174) );
  NAND4X1 U271 ( .A(n438), .B(n419), .C(n437), .D(n418), .Y(n169) );
  AND2X1 U272 ( .A(norm_reg[15]), .B(n30), .Y(arg_a[17]) );
  OAI22X1 U273 ( .A(md4[1]), .B(n27), .C(n439), .D(n199), .Y(arg_b[2]) );
  OAI22X1 U274 ( .A(n31), .B(n130), .C(n146), .D(n33), .Y(arg_a[2]) );
  OAI22X1 U275 ( .A(md4[2]), .B(n27), .C(n147), .D(n199), .Y(arg_b[3]) );
  OAI22X1 U276 ( .A(n30), .B(n140), .C(n425), .D(n33), .Y(arg_a[3]) );
  OAI22X1 U277 ( .A(md4[3]), .B(n27), .C(n438), .D(n199), .Y(arg_b[4]) );
  OAI22X1 U278 ( .A(n30), .B(n131), .C(n154), .D(n33), .Y(arg_a[4]) );
  OAI22X1 U279 ( .A(md4[2]), .B(n26), .C(n193), .D(n147), .Y(arg_d[3]) );
  OAI222XL U280 ( .A(n12), .B(n94), .C(n195), .D(n146), .E(n32), .F(n91), .Y(
        arg_c[3]) );
  OAI22X1 U281 ( .A(md4[4]), .B(n27), .C(n419), .D(n199), .Y(arg_b[5]) );
  OAI22X1 U282 ( .A(n30), .B(n141), .C(n426), .D(n33), .Y(arg_a[5]) );
  OAI22X1 U283 ( .A(md4[3]), .B(n26), .C(n193), .D(n438), .Y(arg_d[4]) );
  OAI222XL U284 ( .A(n194), .B(n92), .C(n7), .D(n425), .E(arg_a[0]), .F(n90), 
        .Y(arg_c[4]) );
  OAI22X1 U285 ( .A(md4[5]), .B(n27), .C(n437), .D(n199), .Y(arg_b[6]) );
  OAI22X1 U286 ( .A(n30), .B(n132), .C(n155), .D(n34), .Y(arg_a[6]) );
  OAI22X1 U287 ( .A(md4[4]), .B(n26), .C(n193), .D(n419), .Y(arg_d[5]) );
  OAI222XL U288 ( .A(n12), .B(n91), .C(n195), .D(n154), .E(arg_a[0]), .F(n89), 
        .Y(arg_c[5]) );
  OAI22X1 U289 ( .A(md4[6]), .B(n27), .C(n418), .D(n199), .Y(arg_b[7]) );
  OAI22X1 U290 ( .A(n30), .B(n142), .C(n427), .D(n34), .Y(arg_a[7]) );
  OAI22X1 U291 ( .A(md4[5]), .B(n26), .C(n193), .D(n437), .Y(arg_d[6]) );
  OAI222XL U292 ( .A(n194), .B(n90), .C(n7), .D(n426), .E(arg_a[0]), .F(n88), 
        .Y(arg_c[6]) );
  OAI22X1 U293 ( .A(md4[7]), .B(n28), .C(n436), .D(n199), .Y(arg_b[8]) );
  OAI22X1 U294 ( .A(n30), .B(n133), .C(n156), .D(n33), .Y(arg_a[8]) );
  OAI22X1 U295 ( .A(md4[6]), .B(n26), .C(n193), .D(n418), .Y(arg_d[7]) );
  OAI222XL U296 ( .A(n12), .B(n89), .C(n195), .D(n155), .E(n32), .F(n87), .Y(
        arg_c[7]) );
  OAI22X1 U297 ( .A(md5[0]), .B(n192), .C(n417), .D(n199), .Y(arg_b[9]) );
  OAI22X1 U298 ( .A(n30), .B(n143), .C(n428), .D(n34), .Y(arg_a[9]) );
  OAI22X1 U299 ( .A(md4[7]), .B(n26), .C(n193), .D(n436), .Y(arg_d[8]) );
  OAI222XL U300 ( .A(n194), .B(n88), .C(n7), .D(n427), .E(n32), .F(n86), .Y(
        arg_c[8]) );
  OAI22X1 U301 ( .A(md5[1]), .B(n28), .C(n435), .D(n13), .Y(arg_b[10]) );
  OAI22X1 U302 ( .A(n30), .B(n134), .C(n157), .D(n34), .Y(arg_a[10]) );
  OAI22X1 U303 ( .A(md5[0]), .B(n192), .C(n193), .D(n417), .Y(arg_d[9]) );
  OAI222XL U304 ( .A(n12), .B(n87), .C(n195), .D(n156), .E(n31), .F(n85), .Y(
        arg_c[9]) );
  OAI22X1 U305 ( .A(md5[2]), .B(n28), .C(n416), .D(n13), .Y(arg_b[11]) );
  OAI22X1 U306 ( .A(n31), .B(n144), .C(n429), .D(n34), .Y(arg_a[11]) );
  OAI22X1 U307 ( .A(md5[1]), .B(n192), .C(n17), .D(n435), .Y(arg_d[10]) );
  OAI222XL U308 ( .A(n194), .B(n86), .C(n7), .D(n428), .E(n31), .F(n84), .Y(
        arg_c[10]) );
  OAI22X1 U309 ( .A(md5[3]), .B(n28), .C(n434), .D(n13), .Y(arg_b[12]) );
  OAI22X1 U310 ( .A(n31), .B(n135), .C(n158), .D(n33), .Y(arg_a[12]) );
  OAI22X1 U311 ( .A(md5[2]), .B(n192), .C(n17), .D(n416), .Y(arg_d[11]) );
  OAI222XL U312 ( .A(n12), .B(n85), .C(n195), .D(n157), .E(n31), .F(n83), .Y(
        arg_c[11]) );
  OAI22X1 U313 ( .A(md5[4]), .B(n28), .C(n415), .D(n13), .Y(arg_b[13]) );
  OAI22X1 U314 ( .A(n31), .B(n145), .C(n430), .D(n34), .Y(arg_a[13]) );
  OAI22X1 U315 ( .A(md5[3]), .B(n192), .C(n17), .D(n434), .Y(arg_d[12]) );
  OAI222XL U316 ( .A(n194), .B(n84), .C(n7), .D(n429), .E(arg_a[0]), .F(n82), 
        .Y(arg_c[12]) );
  OAI22X1 U317 ( .A(md5[5]), .B(n27), .C(n433), .D(n13), .Y(arg_b[14]) );
  OAI22X1 U318 ( .A(n31), .B(n136), .C(n159), .D(n34), .Y(arg_a[14]) );
  OAI22X1 U319 ( .A(md5[4]), .B(n192), .C(n17), .D(n415), .Y(arg_d[13]) );
  OAI222XL U320 ( .A(n12), .B(n83), .C(n195), .D(n158), .E(arg_a[0]), .F(n81), 
        .Y(arg_c[13]) );
  OAI22X1 U321 ( .A(md5[6]), .B(n27), .C(n160), .D(n13), .Y(arg_b[15]) );
  OAI22X1 U322 ( .A(n31), .B(n137), .C(n431), .D(n34), .Y(arg_a[15]) );
  OAI22X1 U323 ( .A(md5[5]), .B(n192), .C(n17), .D(n433), .Y(arg_d[14]) );
  OAI222XL U324 ( .A(n194), .B(n82), .C(n7), .D(n430), .E(n32), .F(n80), .Y(
        arg_c[14]) );
  OAI22X1 U325 ( .A(md5[6]), .B(n192), .C(n17), .D(n160), .Y(arg_d[15]) );
  OAI222XL U326 ( .A(n12), .B(n81), .C(n195), .D(n159), .E(n32), .F(n79), .Y(
        arg_c[15]) );
  INVX1 U327 ( .A(sum1[16]), .Y(n79) );
  OAI22X1 U328 ( .A(md4[1]), .B(n26), .C(n193), .D(n439), .Y(arg_d[2]) );
  OAI222XL U329 ( .A(n194), .B(n95), .C(sum1[17]), .D(n196), .E(n32), .F(n92), 
        .Y(arg_c[2]) );
  INVX1 U330 ( .A(sum1[1]), .Y(n95) );
  OAI22X1 U331 ( .A(md5[7]), .B(n27), .C(n432), .D(n13), .Y(arg_b[16]) );
  ENOX1 U332 ( .A(n32), .B(n148), .C(norm_reg[14]), .D(n32), .Y(arg_a[16]) );
  OAI22X1 U333 ( .A(md5[7]), .B(n28), .C(n17), .D(n432), .Y(arg_d[16]) );
  OAI222XL U334 ( .A(n194), .B(n80), .C(n7), .D(n431), .E(n32), .F(n68), .Y(
        arg_c[16]) );
  AOI21X1 U335 ( .B(mdu_op[0]), .C(mdu_op[1]), .A(n28), .Y(arg_a[0]) );
  NOR21XL U336 ( .B(arg_c[0]), .A(n198), .Y(arg_c[17]) );
  AOI22X1 U337 ( .A(norm_reg[14]), .B(n68), .C(sum1[16]), .D(sum1[17]), .Y(
        n198) );
  OAI22X1 U338 ( .A(md4[0]), .B(n27), .C(n153), .D(n199), .Y(arg_b[1]) );
  OAI21X1 U339 ( .B(n32), .C(n139), .A(n196), .Y(arg_a[1]) );
  OAI22X1 U340 ( .A(n185), .B(n39), .C(n268), .D(n275), .Y(N485) );
  AOI222XL U341 ( .A(sum[10]), .B(n22), .C(n18), .D(norm_reg[7]), .E(n262), 
        .F(sum1[9]), .Y(n275) );
  OAI22X1 U342 ( .A(n5), .B(n41), .C(n268), .D(n273), .Y(N487) );
  AOI222XL U343 ( .A(sum[12]), .B(n21), .C(n259), .D(norm_reg[9]), .E(n262), 
        .F(sum1[11]), .Y(n273) );
  OAI22X1 U344 ( .A(n43), .B(n5), .C(n268), .D(n271), .Y(N489) );
  AOI222XL U345 ( .A(sum[14]), .B(n21), .C(n259), .D(norm_reg[11]), .E(n262), 
        .F(sum1[13]), .Y(n271) );
  OAI22X1 U346 ( .A(n185), .B(n45), .C(n268), .D(n269), .Y(N491) );
  AOI222XL U347 ( .A(sum[16]), .B(n22), .C(n18), .D(norm_reg[13]), .E(n262), 
        .F(sum1[15]), .Y(n269) );
  OAI22X1 U348 ( .A(n5), .B(n38), .C(n268), .D(n276), .Y(N484) );
  AOI222XL U349 ( .A(sum[9]), .B(n21), .C(n259), .D(norm_reg[6]), .E(n262), 
        .F(sum1[8]), .Y(n276) );
  OAI22X1 U350 ( .A(n185), .B(n40), .C(n268), .D(n274), .Y(N486) );
  AOI222XL U351 ( .A(sum[11]), .B(n22), .C(n18), .D(norm_reg[8]), .E(n262), 
        .F(sum1[10]), .Y(n274) );
  OAI22X1 U352 ( .A(n5), .B(n42), .C(n268), .D(n272), .Y(N488) );
  AOI222XL U353 ( .A(sum[13]), .B(n21), .C(n259), .D(norm_reg[10]), .E(n262), 
        .F(sum1[12]), .Y(n272) );
  OAI22X1 U354 ( .A(n185), .B(n44), .C(n268), .D(n270), .Y(N490) );
  AOI222XL U355 ( .A(sum[15]), .B(n22), .C(n18), .D(norm_reg[12]), .E(n262), 
        .F(sum1[14]), .Y(n270) );
  OAI22X1 U356 ( .A(n191), .B(n41), .C(n283), .D(n69), .Y(N457) );
  AOI222XL U357 ( .A(sum[4]), .B(n22), .C(n259), .D(norm_reg[1]), .E(n14), .F(
        sum1[3]), .Y(n283) );
  OAI22X1 U358 ( .A(n43), .B(n191), .C(n281), .D(n69), .Y(N459) );
  AOI222XL U359 ( .A(sum[6]), .B(n22), .C(n259), .D(norm_reg[3]), .E(n14), .F(
        sum1[5]), .Y(n281) );
  OAI22X1 U360 ( .A(n191), .B(n45), .C(n279), .D(n69), .Y(N461) );
  AOI222XL U361 ( .A(sum[8]), .B(n21), .C(n18), .D(norm_reg[5]), .E(n14), .F(
        sum1[7]), .Y(n279) );
  OAI22X1 U362 ( .A(n191), .B(n42), .C(n282), .D(n69), .Y(N458) );
  AOI222XL U363 ( .A(sum[5]), .B(n21), .C(n18), .D(norm_reg[2]), .E(n14), .F(
        sum1[4]), .Y(n282) );
  OAI22X1 U364 ( .A(n191), .B(n44), .C(n280), .D(n69), .Y(N460) );
  AOI222XL U365 ( .A(sum[7]), .B(n22), .C(n259), .D(norm_reg[4]), .E(n14), .F(
        sum1[6]), .Y(n280) );
  OAI22X1 U366 ( .A(n191), .B(n40), .C(n284), .D(n69), .Y(N456) );
  AOI222XL U367 ( .A(sum[3]), .B(n22), .C(n18), .D(norm_reg[0]), .E(n14), .F(
        sum1[2]), .Y(n284) );
  NOR2X1 U368 ( .A(mdu_op[0]), .B(mdu_op[1]), .Y(n192) );
  NAND2X1 U369 ( .A(md0[0]), .B(n26), .Y(n199) );
  OAI32X1 U370 ( .A(n264), .B(n265), .C(n266), .D(n8), .E(n93), .Y(N566) );
  AOI22X1 U371 ( .A(n109), .B(md3[6]), .C(md1[6]), .D(n263), .Y(n266) );
  INVX1 U372 ( .A(sum[1]), .Y(n93) );
  OAI22X1 U373 ( .A(n44), .B(n186), .C(n292), .D(n298), .Y(N412) );
  AOI221XL U374 ( .A(n299), .B(md3[7]), .C(md3[5]), .D(n300), .E(n301), .Y(
        n298) );
  OAI22X1 U375 ( .A(n54), .B(n302), .C(n303), .D(n145), .Y(n301) );
  OAI22X1 U376 ( .A(n45), .B(n186), .C(n292), .D(n293), .Y(N413) );
  AOI221XL U377 ( .A(md3[5]), .B(n294), .C(n16), .D(n21), .E(n295), .Y(n293)
         );
  OAI22X1 U378 ( .A(n178), .B(n296), .C(n137), .D(n297), .Y(n295) );
  OAI22X1 U379 ( .A(n38), .B(n367), .C(n368), .D(n385), .Y(N191) );
  AOI222XL U380 ( .A(n382), .B(n21), .C(n299), .D(md0[1]), .E(md0[2]), .F(n384), .Y(n385) );
  NOR2X1 U381 ( .A(n97), .B(mdu_op[0]), .Y(n200) );
  EORX1 U382 ( .A(n200), .B(md3[7]), .C(n197), .D(n129), .Y(n196) );
  OAI22X1 U383 ( .A(n42), .B(n186), .C(n292), .D(n307), .Y(N410) );
  AOI221XL U384 ( .A(md3[2]), .B(n99), .C(n102), .D(sum[14]), .E(n308), .Y(
        n307) );
  OAI222XL U385 ( .A(n136), .B(n24), .C(n137), .D(n306), .E(n104), .F(n135), 
        .Y(n308) );
  OAI22X1 U386 ( .A(n43), .B(n186), .C(n292), .D(n304), .Y(N411) );
  AOI221XL U387 ( .A(md3[3]), .B(n99), .C(n102), .D(sum[15]), .E(n305), .Y(
        n304) );
  OAI222XL U388 ( .A(n137), .B(n25), .C(n148), .D(n306), .E(n104), .F(n145), 
        .Y(n305) );
  NAND2X1 U389 ( .A(mdu_op[0]), .B(n97), .Y(n197) );
  INVX1 U390 ( .A(mdu_op[1]), .Y(n97) );
  INVX1 U391 ( .A(md1[7]), .Y(n129) );
  OAI22X1 U392 ( .A(n41), .B(n186), .C(n292), .D(n309), .Y(N409) );
  AOI221XL U393 ( .A(md3[1]), .B(n99), .C(n102), .D(sum[13]), .E(n310), .Y(
        n309) );
  OAI222XL U394 ( .A(n145), .B(n24), .C(n136), .D(n306), .E(n104), .F(n144), 
        .Y(n310) );
  INVX1 U395 ( .A(md2[1]), .Y(n130) );
  INVX1 U396 ( .A(md2[0]), .Y(n139) );
  INVX1 U397 ( .A(md4[1]), .Y(n439) );
  INVX1 U398 ( .A(md4[0]), .Y(n153) );
  INVX1 U399 ( .A(norm_reg[0]), .Y(n146) );
  OAI22X1 U400 ( .A(n40), .B(n186), .C(n292), .D(n311), .Y(N408) );
  AOI221XL U401 ( .A(md3[0]), .B(n99), .C(n102), .D(sum[12]), .E(n312), .Y(
        n311) );
  OAI222XL U402 ( .A(n135), .B(n24), .C(n145), .D(n306), .E(n104), .F(n134), 
        .Y(n312) );
  OAI22X1 U403 ( .A(n39), .B(n186), .C(n292), .D(n313), .Y(N407) );
  AOI221XL U404 ( .A(md2[7]), .B(n99), .C(n102), .D(sum[11]), .E(n314), .Y(
        n313) );
  OAI222XL U405 ( .A(n144), .B(n24), .C(n135), .D(n306), .E(n104), .F(n143), 
        .Y(n314) );
  INVX1 U406 ( .A(md4[2]), .Y(n147) );
  INVX1 U407 ( .A(md2[2]), .Y(n140) );
  INVX1 U408 ( .A(norm_reg[1]), .Y(n425) );
  OAI22X1 U409 ( .A(n38), .B(n186), .C(n292), .D(n315), .Y(N406) );
  AOI221XL U410 ( .A(md2[6]), .B(n99), .C(n102), .D(sum[10]), .E(n316), .Y(
        n315) );
  OAI222XL U411 ( .A(n134), .B(n24), .C(n144), .D(n306), .E(n104), .F(n133), 
        .Y(n316) );
  INVX1 U412 ( .A(md2[3]), .Y(n131) );
  INVX1 U413 ( .A(md2[4]), .Y(n141) );
  INVX1 U414 ( .A(md4[4]), .Y(n419) );
  INVX1 U415 ( .A(md4[3]), .Y(n438) );
  INVX1 U416 ( .A(norm_reg[2]), .Y(n154) );
  INVX1 U417 ( .A(norm_reg[3]), .Y(n426) );
  OAI22X1 U418 ( .A(n45), .B(n187), .C(n319), .D(n320), .Y(N340) );
  AOI221XL U419 ( .A(md2[5]), .B(n99), .C(n102), .D(sum[9]), .E(n321), .Y(n320) );
  OAI222XL U420 ( .A(n143), .B(n24), .C(n134), .D(n20), .E(n104), .F(n142), 
        .Y(n321) );
  INVX1 U421 ( .A(md4[5]), .Y(n437) );
  INVX1 U422 ( .A(md2[5]), .Y(n132) );
  INVX1 U423 ( .A(norm_reg[4]), .Y(n155) );
  OAI22X1 U424 ( .A(n44), .B(n187), .C(n319), .D(n322), .Y(N339) );
  AOI221XL U425 ( .A(md2[4]), .B(n99), .C(n102), .D(sum[8]), .E(n323), .Y(n322) );
  OAI222XL U426 ( .A(n133), .B(n24), .C(n143), .D(n20), .E(n11), .F(n132), .Y(
        n323) );
  OAI22X1 U427 ( .A(n43), .B(n187), .C(n319), .D(n324), .Y(N338) );
  AOI221XL U428 ( .A(md2[3]), .B(n99), .C(n102), .D(sum[7]), .E(n325), .Y(n324) );
  OAI222XL U429 ( .A(n142), .B(n24), .C(n133), .D(n20), .E(n11), .F(n141), .Y(
        n325) );
  INVX1 U430 ( .A(md4[6]), .Y(n418) );
  INVX1 U431 ( .A(md2[7]), .Y(n133) );
  INVX1 U432 ( .A(md2[6]), .Y(n142) );
  INVX1 U433 ( .A(md4[7]), .Y(n436) );
  INVX1 U434 ( .A(norm_reg[5]), .Y(n427) );
  INVX1 U435 ( .A(norm_reg[6]), .Y(n156) );
  NAND3X1 U436 ( .A(n186), .B(n187), .C(n188), .Y(n413) );
  NAND31X1 U437 ( .C(n189), .A(n46), .B(set_div32), .Y(n188) );
  OAI22X1 U438 ( .A(n40), .B(n187), .C(n319), .D(n330), .Y(N335) );
  AOI221XL U439 ( .A(md2[0]), .B(n99), .C(n102), .D(sum[4]), .E(n331), .Y(n330) );
  OAI222XL U440 ( .A(n131), .B(n101), .C(n141), .D(n20), .E(n104), .F(n130), 
        .Y(n331) );
  OAI22X1 U441 ( .A(n38), .B(n187), .C(n319), .D(n334), .Y(N333) );
  AOI221XL U442 ( .A(md1[6]), .B(n6), .C(n16), .D(sum[2]), .E(n335), .Y(n334)
         );
  OAI222XL U443 ( .A(n130), .B(n101), .C(n140), .D(n20), .E(n104), .F(n129), 
        .Y(n335) );
  OAI22X1 U444 ( .A(n44), .B(n345), .C(n190), .D(n349), .Y(N265) );
  AOI221XL U445 ( .A(md1[4]), .B(n15), .C(n341), .D(sum1[1]), .E(n350), .Y(
        n349) );
  OAI222XL U446 ( .A(n129), .B(n101), .C(n139), .D(n306), .E(n106), .F(n128), 
        .Y(n350) );
  OAI22X1 U447 ( .A(n41), .B(n187), .C(n319), .D(n328), .Y(N336) );
  AOI221XL U448 ( .A(md2[1]), .B(n6), .C(n16), .D(sum[5]), .E(n329), .Y(n328)
         );
  OAI222XL U449 ( .A(n141), .B(n101), .C(n132), .D(n20), .E(n11), .F(n140), 
        .Y(n329) );
  OAI22X1 U450 ( .A(n39), .B(n187), .C(n319), .D(n332), .Y(N334) );
  AOI221XL U451 ( .A(md1[7]), .B(n6), .C(n16), .D(sum[3]), .E(n333), .Y(n332)
         );
  OAI222XL U452 ( .A(n140), .B(n101), .C(n131), .D(n20), .E(n104), .F(n139), 
        .Y(n333) );
  OAI22X1 U453 ( .A(n45), .B(n345), .C(n190), .D(n346), .Y(N266) );
  AOI221XL U454 ( .A(md1[5]), .B(n15), .C(n341), .D(sum[1]), .E(n348), .Y(n346) );
  OAI222XL U455 ( .A(n139), .B(n101), .C(n130), .D(n306), .E(n106), .F(n138), 
        .Y(n348) );
  OAI22X1 U456 ( .A(n43), .B(n345), .C(n190), .D(n352), .Y(N264) );
  AOI221XL U457 ( .A(md1[4]), .B(n351), .C(md1[3]), .D(n347), .E(n353), .Y(
        n352) );
  OAI22X1 U458 ( .A(n100), .B(n129), .C(n138), .D(n25), .Y(n353) );
  OAI22X1 U459 ( .A(n42), .B(n345), .C(n190), .D(n354), .Y(N263) );
  AOI221XL U460 ( .A(md1[3]), .B(n351), .C(md1[2]), .D(n347), .E(n355), .Y(
        n354) );
  OAI22X1 U461 ( .A(n100), .B(n138), .C(n101), .D(n128), .Y(n355) );
  OAI22X1 U462 ( .A(n41), .B(n345), .C(n190), .D(n356), .Y(N262) );
  AOI221XL U463 ( .A(md1[2]), .B(n351), .C(md1[1]), .D(n347), .E(n357), .Y(
        n356) );
  OAI22X1 U464 ( .A(n100), .B(n128), .C(n101), .D(n127), .Y(n357) );
  OAI22X1 U465 ( .A(n40), .B(n345), .C(n190), .D(n358), .Y(N261) );
  AOI221XL U466 ( .A(md1[1]), .B(n351), .C(md1[0]), .D(n347), .E(n359), .Y(
        n358) );
  OAI22X1 U467 ( .A(n100), .B(n127), .C(n101), .D(n126), .Y(n359) );
  OAI22X1 U468 ( .A(n39), .B(n345), .C(n190), .D(n360), .Y(N260) );
  AOI221XL U469 ( .A(md1[0]), .B(n351), .C(md0[7]), .D(n347), .E(n361), .Y(
        n360) );
  OAI22X1 U470 ( .A(n100), .B(n126), .C(n25), .D(n125), .Y(n361) );
  OAI22X1 U471 ( .A(n38), .B(n345), .C(n190), .D(n362), .Y(N259) );
  AOI221XL U472 ( .A(md0[7]), .B(n351), .C(md0[6]), .D(n347), .E(n363), .Y(
        n362) );
  OAI22X1 U473 ( .A(n100), .B(n125), .C(n25), .D(n124), .Y(n363) );
  OAI22X1 U474 ( .A(n45), .B(n367), .C(n368), .D(n369), .Y(N198) );
  AOI221XL U475 ( .A(md0[6]), .B(n351), .C(md0[5]), .D(n347), .E(n370), .Y(
        n369) );
  OAI22X1 U476 ( .A(n100), .B(n124), .C(n25), .D(n123), .Y(n370) );
  OAI22X1 U477 ( .A(n44), .B(n367), .C(n368), .D(n371), .Y(N197) );
  AOI221XL U478 ( .A(md0[5]), .B(n351), .C(md0[4]), .D(n347), .E(n372), .Y(
        n371) );
  OAI22X1 U479 ( .A(n100), .B(n123), .C(n25), .D(n122), .Y(n372) );
  OAI22X1 U480 ( .A(n43), .B(n367), .C(n368), .D(n373), .Y(N196) );
  AOI221XL U481 ( .A(md0[4]), .B(n351), .C(md0[3]), .D(n347), .E(n374), .Y(
        n373) );
  OAI22X1 U482 ( .A(n100), .B(n122), .C(n25), .D(n121), .Y(n374) );
  OAI22X1 U483 ( .A(n42), .B(n367), .C(n368), .D(n375), .Y(N195) );
  AOI221XL U484 ( .A(md0[3]), .B(n10), .C(md0[2]), .D(n15), .E(n376), .Y(n375)
         );
  OAI22X1 U485 ( .A(n100), .B(n121), .C(n25), .D(n120), .Y(n376) );
  OAI22X1 U486 ( .A(n41), .B(n367), .C(n368), .D(n377), .Y(N194) );
  AOI221XL U487 ( .A(md0[2]), .B(n10), .C(md0[1]), .D(n15), .E(n378), .Y(n377)
         );
  OAI22X1 U488 ( .A(n4), .B(n120), .C(n25), .D(n119), .Y(n378) );
  OAI22X1 U489 ( .A(n40), .B(n367), .C(n368), .D(n379), .Y(N193) );
  AOI221XL U490 ( .A(md0[1]), .B(n10), .C(md0[0]), .D(n15), .E(n380), .Y(n379)
         );
  OAI22X1 U491 ( .A(n4), .B(n119), .C(n25), .D(n118), .Y(n380) );
  OAI22X1 U492 ( .A(n39), .B(n367), .C(n368), .D(n381), .Y(N192) );
  AOI221XL U493 ( .A(md0[0]), .B(n10), .C(n382), .D(sum1[17]), .E(n383), .Y(
        n381) );
  ENOX1 U494 ( .A(n4), .B(n118), .C(n299), .D(md0[2]), .Y(n383) );
  OAI22X1 U495 ( .A(n42), .B(n187), .C(n319), .D(n326), .Y(N337) );
  AOI221XL U496 ( .A(md2[2]), .B(n6), .C(n16), .D(sum[6]), .E(n327), .Y(n326)
         );
  OAI222XL U497 ( .A(n132), .B(n24), .C(n142), .D(n20), .E(n11), .F(n131), .Y(
        n327) );
  OAI21BX1 U498 ( .C(set_div16), .B(n190), .A(n191), .Y(n414) );
  OAI2B11X1 U499 ( .D(mdu_op[0]), .C(n183), .A(n184), .B(n71), .Y(n411) );
  NAND31X1 U500 ( .C(n5), .A(n78), .B(set_div16), .Y(n184) );
  AOI21X1 U501 ( .B(n221), .C(n222), .A(n201), .Y(N893) );
  NOR32XL U502 ( .B(n223), .C(n212), .A(n224), .Y(n222) );
  AOI211X1 U503 ( .C(n115), .D(n213), .A(n225), .B(n226), .Y(n221) );
  OAI22X1 U504 ( .A(n197), .B(n208), .C(arcon[5]), .D(n219), .Y(n224) );
  INVX1 U505 ( .A(md3[0]), .Y(n143) );
  OAI211X1 U506 ( .C(n201), .D(n215), .A(n5), .B(n71), .Y(N894) );
  AOI211X1 U507 ( .C(n113), .D(n148), .A(n216), .B(n217), .Y(n215) );
  OAI22AX1 U508 ( .D(n209), .C(n210), .A(mdu_op[0]), .B(n208), .Y(n217) );
  OAI221X1 U509 ( .A(n112), .B(n218), .C(n167), .D(n203), .E(n219), .Y(n216)
         );
  INVX1 U510 ( .A(md5[0]), .Y(n417) );
  INVX1 U511 ( .A(norm_reg[7]), .Y(n428) );
  OAI22X1 U512 ( .A(md4[0]), .B(n26), .C(n193), .D(n153), .Y(arg_d[1]) );
  OAI222XL U513 ( .A(n96), .B(n137), .C(n31), .D(n94), .E(n197), .F(n138), .Y(
        arg_c[1]) );
  INVX1 U514 ( .A(md3[2]), .Y(n144) );
  INVX1 U515 ( .A(md5[2]), .Y(n416) );
  INVX1 U516 ( .A(md3[1]), .Y(n134) );
  INVX1 U517 ( .A(md5[1]), .Y(n435) );
  INVX1 U518 ( .A(norm_reg[8]), .Y(n157) );
  INVX1 U519 ( .A(norm_reg[9]), .Y(n429) );
  INVX1 U520 ( .A(md3[3]), .Y(n135) );
  INVX1 U521 ( .A(md5[3]), .Y(n434) );
  INVX1 U522 ( .A(norm_reg[10]), .Y(n158) );
  INVX1 U523 ( .A(md3[4]), .Y(n145) );
  INVX1 U524 ( .A(md5[4]), .Y(n415) );
  INVX1 U525 ( .A(md3[5]), .Y(n136) );
  NAND2X1 U526 ( .A(n180), .B(n181), .Y(n410) );
  NAND3X1 U527 ( .A(n182), .B(n47), .C(setmdef), .Y(n180) );
  NAND3X1 U528 ( .A(n182), .B(n46), .C(arcon[7]), .Y(n181) );
  NAND2X1 U529 ( .A(sfroe), .B(n72), .Y(n182) );
  INVX1 U530 ( .A(md5[5]), .Y(n433) );
  INVX1 U531 ( .A(norm_reg[11]), .Y(n430) );
  INVX1 U532 ( .A(norm_reg[12]), .Y(n159) );
  INVX1 U533 ( .A(md3[6]), .Y(n137) );
  INVX1 U534 ( .A(md5[6]), .Y(n160) );
  INVX1 U535 ( .A(norm_reg[13]), .Y(n431) );
  NAND2X1 U536 ( .A(md0[1]), .B(n26), .Y(n193) );
  INVX1 U537 ( .A(md3[7]), .Y(n148) );
  INVX1 U538 ( .A(md5[7]), .Y(n432) );
  INVX1 U539 ( .A(md1[6]), .Y(n138) );
  AOI21BBXL U540 ( .B(md3[6]), .C(n296), .A(n294), .Y(n303) );
  AOI222XL U541 ( .A(N613), .B(n392), .C(N97), .D(n393), .E(arcon[3]), .F(n394), .Y(n249) );
  AOI222XL U542 ( .A(N614), .B(n392), .C(N98), .D(n393), .E(arcon[4]), .F(n394), .Y(n247) );
  AOI222XL U543 ( .A(N612), .B(n392), .C(N96), .D(n393), .E(arcon[2]), .F(n394), .Y(n250) );
  AOI222XL U544 ( .A(n420), .B(n392), .C(N95), .D(n393), .E(arcon[1]), .F(n394), .Y(n251) );
  AOI222XL U545 ( .A(N610), .B(n392), .C(n150), .D(n393), .E(arcon[0]), .F(
        n394), .Y(n252) );
  NOR2X1 U546 ( .A(oper_reg[3]), .B(oper_reg[2]), .Y(n399) );
  NOR2X1 U547 ( .A(oper_reg[1]), .B(oper_reg[0]), .Y(n405) );
  NOR2X1 U548 ( .A(n114), .B(oper_reg[1]), .Y(n389) );
  NOR2X1 U549 ( .A(n152), .B(oper_reg[2]), .Y(n402) );
  NAND3X1 U550 ( .A(n405), .B(oper_reg[3]), .C(oper_reg[2]), .Y(n208) );
  INVX1 U551 ( .A(oper_reg[1]), .Y(n117) );
  INVX1 U552 ( .A(oper_reg[2]), .Y(n149) );
  INVX1 U553 ( .A(oper_reg[3]), .Y(n152) );
  INVX1 U554 ( .A(oper_reg[0]), .Y(n114) );
  OAI221X1 U555 ( .A(md3[6]), .B(n296), .C(n336), .D(n337), .E(n103), .Y(n347)
         );
  NOR2X1 U556 ( .A(n149), .B(oper_reg[3]), .Y(n403) );
  NOR2X1 U557 ( .A(n117), .B(oper_reg[0]), .Y(n400) );
  NAND3X1 U558 ( .A(n389), .B(oper_reg[3]), .C(oper_reg[2]), .Y(n223) );
  NAND43X1 U559 ( .B(arcon[0]), .C(arcon[1]), .D(arcon[2]), .A(n234), .Y(n207)
         );
  NOR2X1 U560 ( .A(arcon[4]), .B(arcon[3]), .Y(n234) );
  OAI31XL U561 ( .A(n206), .B(md3[7]), .C(n207), .D(n167), .Y(n226) );
  NOR4XL U562 ( .A(n422), .B(N610), .C(counter_st[1]), .D(counter_st[3]), .Y(
        n228) );
  NAND2X1 U563 ( .A(counter_st[4]), .B(n228), .Y(n211) );
  INVX1 U564 ( .A(counter_st[4]), .Y(n423) );
  OAI31XL U565 ( .A(n220), .B(N610), .C(n420), .D(n178), .Y(n203) );
  INVX1 U566 ( .A(counter_st[1]), .Y(n420) );
  NAND3X1 U567 ( .A(n424), .B(n423), .C(n422), .Y(n220) );
  INVX1 U568 ( .A(counter_st[2]), .Y(n422) );
  INVX1 U569 ( .A(counter_st[3]), .Y(n424) );
  INVX1 U570 ( .A(N610), .Y(n150) );
  NOR2X1 U571 ( .A(md3[6]), .B(md3[5]), .Y(n178) );
  NAND4X1 U572 ( .A(counter_st[4]), .B(counter_st[1]), .C(n236), .D(n150), .Y(
        n213) );
  NOR2X1 U573 ( .A(counter_st[3]), .B(counter_st[2]), .Y(n236) );
  INVX1 U574 ( .A(md1[5]), .Y(n128) );
  NOR4XL U575 ( .A(md3[7]), .B(md3[4]), .C(md3[3]), .D(md3[2]), .Y(n177) );
  NOR4XL U576 ( .A(md3[1]), .B(md3[0]), .C(md2[7]), .D(md2[6]), .Y(n176) );
  NOR4XL U577 ( .A(md2[5]), .B(md2[4]), .C(md2[3]), .D(md2[2]), .Y(n175) );
  INVX1 U578 ( .A(md1[2]), .Y(n125) );
  NAND4X1 U579 ( .A(n434), .B(n415), .C(n172), .D(n173), .Y(n168) );
  NOR3XL U580 ( .A(md5[5]), .B(md5[7]), .C(md5[6]), .Y(n172) );
  NOR4XL U581 ( .A(md5[2]), .B(md5[1]), .C(md5[0]), .D(md4[7]), .Y(n173) );
  INVX1 U582 ( .A(md0[3]), .Y(n118) );
  INVX1 U583 ( .A(md1[4]), .Y(n127) );
  INVX1 U584 ( .A(md1[3]), .Y(n126) );
  INVX1 U585 ( .A(md1[1]), .Y(n124) );
  INVX1 U586 ( .A(md0[7]), .Y(n122) );
  INVX1 U587 ( .A(md0[6]), .Y(n121) );
  INVX1 U588 ( .A(md0[5]), .Y(n120) );
  INVX1 U589 ( .A(md0[4]), .Y(n119) );
  INVX1 U590 ( .A(md1[0]), .Y(n123) );
  NAND2X1 U591 ( .A(arcon[6]), .B(n167), .Y(n165) );
  INVX1 U592 ( .A(arcon[5]), .Y(n116) );
  INVX1 U593 ( .A(set_div32), .Y(n78) );
  XNOR2XL U594 ( .A(counter_st[4]), .B(r384_carry[4]), .Y(N614) );
  OR2X1 U595 ( .A(r384_carry[3]), .B(counter_st[3]), .Y(r384_carry[4]) );
  XNOR2XL U596 ( .A(r384_carry[3]), .B(counter_st[3]), .Y(N613) );
  OR2X1 U597 ( .A(counter_st[1]), .B(counter_st[2]), .Y(r384_carry[3]) );
  XNOR2XL U598 ( .A(counter_st[1]), .B(counter_st[2]), .Y(N612) );
  OR2X1 U599 ( .A(counter_st[1]), .B(N610), .Y(n49) );
  OAI21BBX1 U600 ( .A(N610), .B(counter_st[1]), .C(n49), .Y(N95) );
  OR2X1 U601 ( .A(n49), .B(counter_st[2]), .Y(n50) );
  OAI21BBX1 U602 ( .A(n49), .B(counter_st[2]), .C(n50), .Y(N96) );
  XNOR2XL U603 ( .A(counter_st[3]), .B(n50), .Y(N97) );
  OR2X1 U604 ( .A(counter_st[3]), .B(n50), .Y(n51) );
  XNOR2XL U605 ( .A(counter_st[4]), .B(n51), .Y(N98) );
endmodule


module mdu_a0_DW01_add_1 ( A, B, CI, SUM, CO );
  input [17:0] A;
  input [17:0] B;
  output [17:0] SUM;
  input CI;
  output CO;

  wire   [17:1] carry;

  FAD1X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .SO(
        SUM[16]) );
  FAD1X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .SO(
        SUM[15]) );
  FAD1X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .SO(
        SUM[14]) );
  FAD1X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .SO(
        SUM[13]) );
  FAD1X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .SO(
        SUM[12]) );
  FAD1X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .SO(
        SUM[11]) );
  FAD1X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .SO(
        SUM[10]) );
  FAD1X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .SO(SUM[9])
         );
  FAD1X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .SO(SUM[8])
         );
  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  XOR2X1 U1 ( .A(A[17]), .B(carry[17]), .Y(SUM[17]) );
  AND2X1 U2 ( .A(B[0]), .B(A[0]), .Y(carry[1]) );
endmodule


module mdu_a0_DW01_add_0 ( A, B, CI, SUM, CO );
  input [17:0] A;
  input [17:0] B;
  output [17:0] SUM;
  input CI;
  output CO;

  wire   [17:1] carry;

  FAD1X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .SO(
        SUM[16]) );
  FAD1X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .SO(
        SUM[15]) );
  FAD1X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .SO(
        SUM[14]) );
  FAD1X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .SO(
        SUM[13]) );
  FAD1X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .SO(
        SUM[12]) );
  FAD1X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .SO(
        SUM[11]) );
  FAD1X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .SO(
        SUM[10]) );
  FAD1X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .SO(SUM[9])
         );
  FAD1X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .SO(SUM[8])
         );
  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  XOR2X1 U1 ( .A(A[17]), .B(carry[17]), .Y(SUM[17]) );
  AND2X1 U2 ( .A(B[0]), .B(A[0]), .Y(carry[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mdu_a0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mdu_a0_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mdu_a0_3 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mdu_a0_4 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mdu_a0_5 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mdu_a0_6 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mdu_a0_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module wakeupctrl_a0 ( irq, int0ff, int1ff, it0, it1, isreg, intprior0, 
        intprior1, eal, eint0, eint1, pmuintreq );
  input [3:0] isreg;
  input [1:0] intprior0;
  input [1:0] intprior1;
  input irq, int0ff, int1ff, it0, it1, eal, eint0, eint1;
  output pmuintreq;
  wire   n6, n7, n8, n9, n10, n11, n12, n1, n2, n3, n4, n5;

  OAI21BX1 U1 ( .C(eal), .B(n6), .A(n1), .Y(pmuintreq) );
  INVX1 U2 ( .A(irq), .Y(n1) );
  AOI33X1 U3 ( .A(eint0), .B(n7), .C(n8), .D(eint1), .E(n9), .F(n10), .Y(n6)
         );
  NOR3XL U4 ( .A(int1ff), .B(it1), .C(isreg[3]), .Y(n10) );
  NOR3XL U5 ( .A(int0ff), .B(it0), .C(isreg[3]), .Y(n8) );
  OAI21X1 U6 ( .B(n3), .C(n5), .A(n12), .Y(n7) );
  GEN2XL U7 ( .D(isreg[0]), .E(n3), .C(isreg[1]), .B(n5), .A(isreg[2]), .Y(n12) );
  INVX1 U8 ( .A(intprior1[0]), .Y(n5) );
  INVX1 U9 ( .A(intprior0[0]), .Y(n3) );
  OAI21X1 U10 ( .B(n2), .C(n4), .A(n11), .Y(n9) );
  GEN2XL U11 ( .D(isreg[0]), .E(n2), .C(isreg[1]), .B(n4), .A(isreg[2]), .Y(
        n11) );
  INVX1 U12 ( .A(intprior1[1]), .Y(n4) );
  INVX1 U13 ( .A(intprior0[1]), .Y(n2) );
endmodule


module pmurstctrl_a0 ( resetff, wdts, srst, pmuintreq, stop, idle, clkcpu_en, 
        clkper_en, cpu_resume, rsttowdt, rsttosrst, rst );
  input resetff, wdts, srst, pmuintreq, stop, idle;
  output clkcpu_en, clkper_en, cpu_resume, rsttowdt, rsttosrst, rst;
  wire   n2;

  OAI21X1 U1 ( .B(stop), .C(idle), .A(n2), .Y(clkcpu_en) );
  NAND2X1 U2 ( .A(stop), .B(n2), .Y(clkper_en) );
  INVX1 U3 ( .A(pmuintreq), .Y(n2) );
  OR2X1 U4 ( .A(srst), .B(resetff), .Y(rsttowdt) );
  OR2X1 U5 ( .A(wdts), .B(rsttowdt), .Y(rst) );
  OR2X1 U6 ( .A(resetff), .B(wdts), .Y(rsttosrst) );
  BUFX3 U7 ( .A(pmuintreq), .Y(cpu_resume) );
endmodule


module sfrmux_a0 ( isfrwait, sfraddr, c, ac, f0, rs, ov, f1, p, acc, b, dpl, 
        dph, dps, dpc, p2, sp, smod, pmw, p2sel, gf0, stop, idle, ckcon, port0, 
        port0ff, rmwinstr, arcon, md0, md1, md2, md3, md4, md5, t0_tmod, 
        t0_tf0, t0_tf1, t0_tr0, t0_tr1, tl0, th0, t1_tmod, t1_tf1, t1_tr1, tl1, 
        th1, wdtrel, ip0wdts, wdt_tm, t2con, s0con, s0buf, s0rell, s0relh, bd, 
        ie0, it0, ie1, it1, iex2, iex3, iex4, iex5, iex6, iex7, iex8, iex9, 
        iex10, iex11, iex12, ien0, ien1, ien2, ip0, ip1, isr_tm, i2c_int, 
        i2cdat_o, i2cadr_o, i2ccon_o, i2csta_o, sfrdatai, tf1_gate, riti0_gate, 
        iex7_gate, iex2_gate, srstflag, int_vect_8b, int_vect_93, int_vect_9b, 
        int_vect_a3, ext_sfr_sel, sfrdatao );
  input [6:0] sfraddr;
  input [1:0] rs;
  input [7:0] acc;
  input [7:0] b;
  input [7:0] dpl;
  input [7:0] dph;
  input [3:0] dps;
  input [5:0] dpc;
  input [7:0] p2;
  input [7:0] sp;
  input [7:0] ckcon;
  input [7:0] port0;
  input [7:0] port0ff;
  input [7:0] arcon;
  input [7:0] md0;
  input [7:0] md1;
  input [7:0] md2;
  input [7:0] md3;
  input [7:0] md4;
  input [7:0] md5;
  input [3:0] t0_tmod;
  input [7:0] tl0;
  input [7:0] th0;
  input [3:0] t1_tmod;
  input [7:0] tl1;
  input [7:0] th1;
  input [7:0] wdtrel;
  input [7:0] t2con;
  input [7:0] s0con;
  input [7:0] s0buf;
  input [7:0] s0rell;
  input [7:0] s0relh;
  input [7:0] ien0;
  input [5:0] ien1;
  input [5:0] ien2;
  input [5:0] ip0;
  input [5:0] ip1;
  input [7:0] i2cdat_o;
  input [7:0] i2cadr_o;
  input [7:0] i2ccon_o;
  input [7:0] i2csta_o;
  input [7:0] sfrdatai;
  output [7:0] sfrdatao;
  input isfrwait, c, ac, f0, ov, f1, p, smod, pmw, p2sel, gf0, stop, idle,
         rmwinstr, t0_tf0, t0_tf1, t0_tr0, t0_tr1, t1_tf1, t1_tr1, ip0wdts,
         wdt_tm, bd, ie0, it0, ie1, it1, iex2, iex3, iex4, iex5, iex6, iex7,
         iex8, iex9, iex10, iex11, iex12, isr_tm, i2c_int, srstflag;
  output tf1_gate, riti0_gate, iex7_gate, iex2_gate, int_vect_8b, int_vect_93,
         int_vect_9b, int_vect_a3, ext_sfr_sel;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347;

  INVXL U2 ( .A(n55), .Y(n64) );
  NAND43X1 U3 ( .B(sfraddr[1]), .C(n25), .D(n28), .A(n70), .Y(n159) );
  NAND21X1 U4 ( .B(n60), .A(n65), .Y(n160) );
  NAND21X1 U5 ( .B(n32), .A(n39), .Y(n60) );
  NAND32XL U6 ( .B(n53), .C(n62), .A(n26), .Y(n148) );
  INVX1 U7 ( .A(n122), .Y(n300) );
  INVX1 U8 ( .A(n52), .Y(n66) );
  NOR3X1 U9 ( .A(n10), .B(n11), .C(n12), .Y(n111) );
  AND2X1 U10 ( .A(sfrdatai[1]), .B(n317), .Y(n12) );
  INVX1 U11 ( .A(n60), .Y(n41) );
  NAND42X1 U12 ( .C(n183), .D(n182), .A(n181), .B(n180), .Y(n184) );
  NOR43XL U13 ( .B(n144), .C(n143), .D(n142), .A(n141), .Y(n185) );
  AOI221XL U14 ( .A(iex7), .B(n252), .C(t2con[0]), .D(n328), .E(n79), .Y(n97)
         );
  INVX1 U15 ( .A(n47), .Y(n337) );
  AOI221XL U16 ( .A(b[7]), .B(n332), .C(arcon[7]), .D(n331), .E(n330), .Y(n333) );
  NAND42X1 U17 ( .C(n288), .D(n287), .A(n286), .B(n285), .Y(sfrdatao[6]) );
  AO2222XL U18 ( .A(md5[6]), .B(n292), .C(md4[6]), .D(n291), .E(md1[6]), .F(
        n290), .G(md3[6]), .H(n289), .Y(n288) );
  AOI221XL U19 ( .A(b[6]), .B(n332), .C(arcon[6]), .D(n331), .E(n284), .Y(n285) );
  AOI221XL U20 ( .A(dpc[4]), .B(n261), .C(ckcon[4]), .D(n298), .E(n238), .Y(
        n244) );
  AOI221XL U21 ( .A(b[4]), .B(n332), .C(arcon[4]), .D(n331), .E(n231), .Y(n248) );
  NAND6XL U22 ( .A(n230), .B(n229), .C(n228), .D(n227), .E(n226), .F(n225), 
        .Y(sfrdatao[3]) );
  AOI221XL U23 ( .A(ien0[3]), .B(n299), .C(ien2[3]), .D(n259), .E(n214), .Y(
        n227) );
  NAND6XL U24 ( .A(n271), .B(n270), .C(n269), .D(n268), .E(n267), .F(n266), 
        .Y(sfrdatao[5]) );
  AOI221XL U25 ( .A(dpc[5]), .B(n261), .C(ckcon[5]), .D(n298), .E(n260), .Y(
        n267) );
  AOI221XL U26 ( .A(b[5]), .B(n332), .C(arcon[5]), .D(n331), .E(n250), .Y(n271) );
  NAND5XL U27 ( .A(n167), .B(n168), .C(n139), .D(n138), .E(n140), .Y(n74) );
  NAND5XL U28 ( .A(n148), .B(n78), .C(n149), .D(n147), .E(n152), .Y(n75) );
  INVX1 U29 ( .A(n51), .Y(n343) );
  NAND6XL U30 ( .A(n129), .B(n118), .C(n133), .D(n128), .E(n130), .F(n50), .Y(
        n51) );
  INVX1 U31 ( .A(n43), .Y(n345) );
  NAND6XL U32 ( .A(n80), .B(n173), .C(n161), .D(n171), .E(n123), .F(n120), .Y(
        n43) );
  NAND2X1 U33 ( .A(s0relh[5]), .B(n318), .Y(n1) );
  NAND2X1 U34 ( .A(port0ff[5]), .B(n341), .Y(n2) );
  NAND2X1 U35 ( .A(sfrdatai[5]), .B(n317), .Y(n3) );
  AND3X1 U36 ( .A(n1), .B(n2), .C(n3), .Y(n256) );
  INVX1 U37 ( .A(n146), .Y(n317) );
  AND2X1 U38 ( .A(s0relh[4]), .B(n318), .Y(n4) );
  AND2X1 U39 ( .A(port0ff[4]), .B(n341), .Y(n5) );
  AND2X2 U40 ( .A(sfrdatai[4]), .B(n317), .Y(n6) );
  NOR3X2 U41 ( .A(n4), .B(n5), .C(n6), .Y(n236) );
  NAND2X1 U42 ( .A(s0relh[3]), .B(n318), .Y(n7) );
  NAND2X1 U43 ( .A(port0ff[3]), .B(n341), .Y(n8) );
  NAND2X1 U44 ( .A(sfrdatai[3]), .B(n317), .Y(n9) );
  AND3X1 U45 ( .A(n7), .B(n8), .C(n9), .Y(n224) );
  NAND32X1 U46 ( .B(n30), .C(n29), .A(n31), .Y(n53) );
  NAND32X2 U47 ( .B(sfraddr[2]), .C(n25), .A(n27), .Y(n71) );
  AND2X1 U48 ( .A(s0relh[1]), .B(n318), .Y(n10) );
  AND2X1 U49 ( .A(port0ff[1]), .B(n341), .Y(n11) );
  NAND21XL U50 ( .B(n60), .A(n64), .Y(n168) );
  NAND32X1 U51 ( .B(sfraddr[5]), .C(n59), .A(n30), .Y(n140) );
  NAND5XL U52 ( .A(sfraddr[3]), .B(sfraddr[6]), .C(n56), .D(n31), .E(n30), .Y(
        n139) );
  AOI221XL U53 ( .A(ien0[1]), .B(n299), .C(ien2[1]), .D(n259), .E(n101), .Y(
        n114) );
  AOI221XL U54 ( .A(iex2), .B(n252), .C(t2con[1]), .D(n328), .E(n103), .Y(n109) );
  NAND21X1 U55 ( .B(sfraddr[6]), .A(n31), .Y(n42) );
  NOR31X1 U56 ( .C(n185), .A(n14), .B(n184), .Y(n210) );
  INVXL U57 ( .A(sfraddr[2]), .Y(n28) );
  NAND21XL U58 ( .B(n67), .A(n65), .Y(n187) );
  NAND21XL U59 ( .B(n69), .A(n68), .Y(n191) );
  NOR5X1 U60 ( .A(n339), .B(n340), .C(n337), .D(n301), .E(n48), .Y(n77) );
  INVX1 U61 ( .A(n46), .Y(n339) );
  INVX1 U62 ( .A(n119), .Y(n340) );
  NAND32XL U63 ( .B(n71), .C(n32), .A(n29), .Y(n59) );
  AOI221XL U64 ( .A(tl1[6]), .B(n306), .C(t1_tmod[2]), .D(n305), .E(n272), .Y(
        n276) );
  INVX2 U65 ( .A(n66), .Y(n17) );
  NAND32X1 U66 ( .B(n31), .C(n29), .A(n30), .Y(n63) );
  NAND32XL U67 ( .B(n29), .C(n42), .A(n30), .Y(n67) );
  INVXL U68 ( .A(n35), .Y(n54) );
  INVXL U69 ( .A(n120), .Y(n261) );
  NAND43X1 U70 ( .B(sfraddr[1]), .C(n67), .D(n28), .A(n25), .Y(n346) );
  INVXL U71 ( .A(n34), .Y(n38) );
  NAND4X1 U72 ( .A(n158), .B(n157), .C(n156), .D(n18), .Y(n14) );
  INVX1 U73 ( .A(n155), .Y(n18) );
  INVX1 U74 ( .A(n210), .Y(n13) );
  AOI221XL U75 ( .A(p2[5]), .B(n311), .C(ien0[5]), .D(n299), .E(n258), .Y(n268) );
  AOI221XL U76 ( .A(p2[4]), .B(n311), .C(ien0[4]), .D(n299), .E(n237), .Y(n245) );
  INVX1 U77 ( .A(n276), .Y(n15) );
  AO222XL U78 ( .A(i2cadr_o[3]), .B(n323), .C(i2cdat_o[3]), .D(n321), .E(rs[0]), .F(n339), .Y(n216) );
  INVX3 U79 ( .A(n194), .Y(n312) );
  INVX3 U80 ( .A(n196), .Y(n295) );
  INVXL U81 ( .A(n161), .Y(n292) );
  INVXL U82 ( .A(n163), .Y(n290) );
  INVX3 U83 ( .A(n193), .Y(n308) );
  INVX3 U84 ( .A(n192), .Y(n309) );
  NAND21XL U85 ( .B(n53), .A(n16), .Y(n129) );
  INVXL U86 ( .A(n78), .Y(n321) );
  INVXL U87 ( .A(n138), .Y(n323) );
  NAND21XL U88 ( .B(n44), .A(n70), .Y(n123) );
  NAND21XL U89 ( .B(n69), .A(n41), .Y(n171) );
  INVXL U90 ( .A(n173), .Y(n332) );
  NAND21XL U91 ( .B(n44), .A(n68), .Y(n198) );
  INVX3 U92 ( .A(n197), .Y(n296) );
  NAND3XL U93 ( .A(n25), .B(n57), .C(n61), .Y(n149) );
  NAND32XL U94 ( .B(n31), .C(n59), .A(n30), .Y(n152) );
  NAND21XL U95 ( .B(n49), .A(n66), .Y(n195) );
  NAND32XL U96 ( .B(sfraddr[6]), .C(n29), .A(n38), .Y(n35) );
  NAND21XL U97 ( .B(n40), .A(n25), .Y(n69) );
  NAND21XL U98 ( .B(n52), .A(n54), .Y(n147) );
  OR2XL U99 ( .A(n25), .B(n40), .Y(n44) );
  NAND21XL U100 ( .B(n67), .A(n64), .Y(n186) );
  INVXL U101 ( .A(n36), .Y(n48) );
  NAND32XL U102 ( .B(n30), .C(n59), .A(n31), .Y(n46) );
  INVXL U103 ( .A(n148), .Y(n322) );
  INVXL U104 ( .A(n133), .Y(n299) );
  NAND32XL U105 ( .B(sfraddr[4]), .C(n42), .A(n29), .Y(n49) );
  NAND32XL U106 ( .B(n63), .C(n62), .A(n26), .Y(n162) );
  NAND32XL U107 ( .B(n26), .C(n63), .A(n61), .Y(n170) );
  NAND32XL U108 ( .B(n27), .C(n26), .A(n28), .Y(n58) );
  NAND32XL U109 ( .B(n33), .C(n28), .A(n27), .Y(n62) );
  NAND32XL U110 ( .B(n53), .C(n55), .A(n32), .Y(n118) );
  NAND21XL U111 ( .B(n55), .A(n54), .Y(n167) );
  NAND21XL U112 ( .B(n31), .A(sfraddr[4]), .Y(n34) );
  INVXL U113 ( .A(sfraddr[6]), .Y(n32) );
  NAND43X1 U114 ( .B(n212), .C(n211), .D(n13), .A(n209), .Y(sfrdatao[2]) );
  NAND42XL U115 ( .C(n316), .D(n315), .A(n314), .B(n313), .Y(n335) );
  NAND43X1 U116 ( .B(n278), .C(n277), .D(n15), .A(n275), .Y(n287) );
  AOI22XL U117 ( .A(acc[7]), .B(n320), .C(i2csta_o[7]), .D(n319), .Y(n326) );
  AOI221X1 U118 ( .A(sfrdatai[6]), .B(n317), .C(port0ff[6]), .D(n341), .E(n279), .Y(n283) );
  NAND6X1 U119 ( .A(n99), .B(n98), .C(n97), .D(n96), .E(n95), .F(n94), .Y(
        sfrdatao[0]) );
  AO222X1 U120 ( .A(th0[6]), .B(n303), .C(md2[6]), .D(n302), .E(th1[6]), .F(
        n301), .Y(n272) );
  AO222XL U121 ( .A(md0[4]), .B(n329), .C(ip1[4]), .D(n249), .E(port0[4]), .F(
        n338), .Y(n231) );
  AO222X1 U122 ( .A(i2cadr_o[1]), .B(n323), .C(i2cdat_o[1]), .D(n321), .E(f1), 
        .F(n339), .Y(n103) );
  NAND21XL U123 ( .B(n36), .A(rmwinstr), .Y(n169) );
  AOI21BXL U124 ( .C(n122), .B(s0con[2]), .A(n121), .Y(n125) );
  AOI21BXL U125 ( .C(n132), .B(ien1[2]), .A(n131), .Y(n135) );
  AOI21BXL U126 ( .C(n173), .B(b[2]), .A(n172), .Y(n174) );
  AO222XL U127 ( .A(md0[6]), .B(n329), .C(t2con[6]), .D(n328), .E(port0[6]), 
        .F(n338), .Y(n284) );
  NAND21XL U128 ( .B(n145), .A(port0ff[2]), .Y(n158) );
  NAND21XL U129 ( .B(n198), .A(wdtrel[2]), .Y(n199) );
  INVXL U130 ( .A(n160), .Y(n302) );
  INVX1 U131 ( .A(n191), .Y(n294) );
  INVX1 U132 ( .A(n187), .Y(n306) );
  INVX1 U133 ( .A(n198), .Y(n293) );
  INVX1 U134 ( .A(n171), .Y(n331) );
  INVX1 U135 ( .A(n123), .Y(n298) );
  INVX1 U136 ( .A(n129), .Y(n259) );
  OR2XL U137 ( .A(n60), .B(n44), .Y(n161) );
  NAND21X1 U138 ( .B(n67), .A(n66), .Y(n196) );
  NAND2X1 U139 ( .A(n41), .B(n66), .Y(n163) );
  NAND21X1 U140 ( .B(n63), .A(n16), .Y(n194) );
  INVX1 U141 ( .A(n67), .Y(n70) );
  INVX1 U142 ( .A(n149), .Y(n319) );
  NOR2X2 U143 ( .A(sfraddr[6]), .B(n17), .Y(n16) );
  INVX1 U144 ( .A(n63), .Y(n39) );
  INVX1 U145 ( .A(n53), .Y(n57) );
  INVX1 U146 ( .A(n168), .Y(n329) );
  INVX1 U147 ( .A(n152), .Y(n320) );
  INVX1 U148 ( .A(n186), .Y(n305) );
  INVX1 U149 ( .A(n195), .Y(n307) );
  INVX1 U150 ( .A(n45), .Y(n347) );
  NAND21X1 U151 ( .B(n300), .A(n198), .Y(n45) );
  INVX1 U152 ( .A(n147), .Y(n318) );
  NAND32XL U153 ( .B(n32), .C(n52), .A(n57), .Y(n78) );
  NAND21X1 U154 ( .B(n59), .A(n38), .Y(n173) );
  NAND32X1 U155 ( .B(n32), .C(n58), .A(n57), .Y(n138) );
  INVXL U156 ( .A(n130), .Y(n311) );
  NAND21X1 U157 ( .B(n58), .A(n68), .Y(n193) );
  NAND21X1 U158 ( .B(n49), .A(n64), .Y(n192) );
  INVX1 U159 ( .A(n49), .Y(n68) );
  INVX1 U160 ( .A(n162), .Y(n289) );
  INVXL U161 ( .A(n159), .Y(n303) );
  INVX1 U162 ( .A(n346), .Y(n301) );
  INVX1 U163 ( .A(n58), .Y(n65) );
  INVX1 U164 ( .A(n62), .Y(n61) );
  INVX1 U165 ( .A(n118), .Y(n297) );
  INVX1 U166 ( .A(n170), .Y(n291) );
  INVX1 U167 ( .A(n128), .Y(n274) );
  INVX1 U168 ( .A(n76), .Y(n342) );
  INVX1 U169 ( .A(n139), .Y(n328) );
  INVX1 U170 ( .A(n145), .Y(n341) );
  INVX1 U171 ( .A(n167), .Y(n249) );
  INVX1 U172 ( .A(n140), .Y(n252) );
  NAND31XL U173 ( .C(n71), .A(n39), .B(n32), .Y(n133) );
  NAND43X1 U174 ( .B(sfraddr[3]), .C(n42), .D(n30), .A(n65), .Y(n120) );
  NAND43XL U175 ( .B(sfraddr[3]), .C(sfraddr[5]), .D(n30), .A(n16), .Y(n119)
         );
  NAND32XL U176 ( .B(n63), .C(n55), .A(n32), .Y(n128) );
  NAND32XL U177 ( .B(n71), .C(n53), .A(n32), .Y(n122) );
  NAND21XL U178 ( .B(n71), .A(n68), .Y(n36) );
  NAND21X1 U179 ( .B(n71), .A(n70), .Y(n197) );
  NAND21XL U180 ( .B(n338), .A(n48), .Y(n145) );
  NAND21X1 U181 ( .B(n28), .A(sfraddr[1]), .Y(n40) );
  NAND32X1 U182 ( .B(n25), .C(n27), .A(n28), .Y(n52) );
  NAND5XL U183 ( .A(sfraddr[6]), .B(sfraddr[5]), .C(sfraddr[4]), .D(n37), .E(
        n29), .Y(n80) );
  INVX1 U184 ( .A(sfraddr[4]), .Y(n30) );
  INVX1 U185 ( .A(n71), .Y(n56) );
  INVX1 U186 ( .A(sfraddr[3]), .Y(n29) );
  INVX3 U187 ( .A(sfraddr[5]), .Y(n31) );
  INVX1 U188 ( .A(sfraddr[1]), .Y(n27) );
  INVX2 U189 ( .A(n26), .Y(n25) );
  NOR21XL U190 ( .B(dps[2]), .A(n119), .Y(n126) );
  NOR5XL U191 ( .A(n341), .B(n340), .C(n339), .D(n338), .E(n337), .Y(n344) );
  NAND42X1 U192 ( .C(n127), .D(n126), .A(n125), .B(n124), .Y(n212) );
  NOR21XL U193 ( .B(n208), .A(n207), .Y(n209) );
  NAND42X1 U194 ( .C(n137), .D(n136), .A(n135), .B(n134), .Y(n211) );
  NAND32XL U195 ( .B(sfraddr[2]), .C(n26), .A(n27), .Y(n55) );
  INVX1 U196 ( .A(n169), .Y(n338) );
  NOR21XL U197 ( .B(p2[2]), .A(n130), .Y(n131) );
  NOR43XL U198 ( .B(n179), .C(n178), .D(n177), .A(n176), .Y(n180) );
  NAND21XL U199 ( .B(n167), .A(ip1[2]), .Y(n179) );
  NAND21X1 U200 ( .B(n175), .A(n174), .Y(n176) );
  NAND21XL U201 ( .B(n168), .A(md0[2]), .Y(n178) );
  AO2222XL U202 ( .A(md5[7]), .B(n292), .C(md4[7]), .D(n291), .E(md1[7]), .F(
        n290), .G(md3[7]), .H(n289), .Y(n336) );
  AO222X1 U203 ( .A(md0[7]), .B(n329), .C(t2con[7]), .D(n328), .E(port0[7]), 
        .F(n338), .Y(n330) );
  AO222XL U204 ( .A(s0buf[3]), .B(n297), .C(s0con[3]), .D(n300), .E(dpc[3]), 
        .F(n261), .Y(n215) );
  AO222XL U205 ( .A(ien1[5]), .B(n257), .C(s0rell[5]), .D(n312), .E(ip0[5]), 
        .F(n274), .Y(n258) );
  AO222X1 U206 ( .A(md5[5]), .B(n292), .C(md4[5]), .D(n291), .E(md3[5]), .F(
        n289), .Y(n251) );
  AO222XL U207 ( .A(s0buf[1]), .B(n297), .C(s0con[1]), .D(n300), .E(dpc[1]), 
        .F(n261), .Y(n102) );
  AO222XL U208 ( .A(ien1[4]), .B(n257), .C(s0rell[4]), .D(n312), .E(ip0[4]), 
        .F(n274), .Y(n237) );
  AO222X1 U209 ( .A(md5[4]), .B(n292), .C(md4[4]), .D(n291), .E(md3[4]), .F(
        n289), .Y(n232) );
  AO2222XL U210 ( .A(s0con[6]), .B(n300), .C(ien0[6]), .D(n299), .E(ckcon[6]), 
        .F(n298), .G(s0buf[6]), .H(n297), .Y(n277) );
  AO2222XL U211 ( .A(s0con[7]), .B(n300), .C(ien0[7]), .D(n299), .E(ckcon[7]), 
        .F(n298), .G(s0buf[7]), .H(n297), .Y(n315) );
  AO2222XL U212 ( .A(wdtrel[6]), .B(n293), .C(tl0[6]), .D(n295), .E(dph[6]), 
        .F(n308), .G(wdt_tm), .H(n294), .Y(n278) );
  AOI22XL U213 ( .A(c), .B(n339), .C(bd), .D(n337), .Y(n324) );
  AOI222XL U214 ( .A(i2cadr_o[7]), .B(n323), .C(i2ccon_o[7]), .D(n322), .E(
        i2cdat_o[7]), .F(n321), .Y(n325) );
  AOI222XL U215 ( .A(wdtrel[3]), .B(n293), .C(tl0[3]), .D(n295), .E(ie1), .F(
        n296), .Y(n229) );
  AOI222XL U216 ( .A(t0_tmod[3]), .B(n305), .C(th1[3]), .D(n301), .E(tl1[3]), 
        .F(n306), .Y(n230) );
  AOI221XL U217 ( .A(ckcon[3]), .B(n298), .C(dps[3]), .D(n340), .E(n215), .Y(
        n226) );
  AND4X1 U218 ( .A(n265), .B(n264), .C(n263), .D(n262), .Y(n266) );
  AOI221XL U219 ( .A(md1[5]), .B(n290), .C(md2[5]), .D(n302), .E(n251), .Y(
        n270) );
  AND4X1 U220 ( .A(n283), .B(n282), .C(n281), .D(n280), .Y(n286) );
  AOI22X1 U221 ( .A(s0relh[6]), .B(n318), .C(acc[6]), .D(n320), .Y(n282) );
  AOI22XL U222 ( .A(i2cadr_o[6]), .B(n323), .C(ac), .D(n339), .Y(n280) );
  AOI222XL U223 ( .A(i2cdat_o[6]), .B(n321), .C(i2csta_o[6]), .D(n319), .E(
        i2ccon_o[6]), .F(n322), .Y(n281) );
  AOI222XL U224 ( .A(i2ccon_o[1]), .B(n322), .C(acc[1]), .D(n320), .E(
        i2csta_o[1]), .F(n319), .Y(n110) );
  AND4X1 U225 ( .A(n107), .B(n106), .C(n105), .D(n104), .Y(n108) );
  AOI222XL U226 ( .A(i2ccon_o[3]), .B(n322), .C(acc[3]), .D(n320), .E(
        i2csta_o[3]), .F(n319), .Y(n223) );
  AND4X1 U227 ( .A(n220), .B(n219), .C(n218), .D(n217), .Y(n221) );
  AOI221X1 U228 ( .A(iex4), .B(n252), .C(t2con[3]), .D(n328), .E(n216), .Y(
        n222) );
  AOI22X1 U229 ( .A(iex5), .B(n252), .C(t2con[4]), .D(n328), .Y(n233) );
  AOI222XL U230 ( .A(rs[1]), .B(n339), .C(i2cdat_o[4]), .D(n321), .E(
        i2cadr_o[4]), .F(n323), .Y(n234) );
  AOI222XL U231 ( .A(i2ccon_o[4]), .B(n322), .C(acc[4]), .D(n320), .E(
        i2csta_o[4]), .F(n319), .Y(n235) );
  AOI22X1 U232 ( .A(iex6), .B(n252), .C(t2con[5]), .D(n328), .Y(n253) );
  AOI222XL U233 ( .A(f0), .B(n339), .C(i2cdat_o[5]), .D(n321), .E(i2cadr_o[5]), 
        .F(n323), .Y(n254) );
  AOI222XL U234 ( .A(i2ccon_o[5]), .B(n322), .C(acc[5]), .D(n320), .E(
        i2csta_o[5]), .F(n319), .Y(n255) );
  AND4X1 U235 ( .A(n242), .B(n241), .C(n240), .D(n239), .Y(n243) );
  AOI221XL U236 ( .A(md1[4]), .B(n290), .C(md2[4]), .D(n302), .E(n232), .Y(
        n247) );
  AOI222XL U237 ( .A(i2ccon_o[0]), .B(n322), .C(acc[0]), .D(n320), .E(
        i2csta_o[0]), .F(n319), .Y(n98) );
  AND4X1 U238 ( .A(n89), .B(n88), .C(n87), .D(n86), .Y(n95) );
  AND4X1 U239 ( .A(n85), .B(n84), .C(n83), .D(n82), .Y(n96) );
  AOI222XL U240 ( .A(wdtrel[1]), .B(n293), .C(tl0[1]), .D(n295), .E(ie0), .F(
        n296), .Y(n116) );
  AOI222XL U241 ( .A(t0_tmod[1]), .B(n305), .C(th1[1]), .D(n301), .E(tl1[1]), 
        .F(n306), .Y(n117) );
  AOI221XL U242 ( .A(ckcon[1]), .B(n298), .C(dps[1]), .D(n340), .E(n102), .Y(
        n113) );
  NAND21XL U243 ( .B(n169), .A(port0[2]), .Y(n177) );
  AND4X1 U244 ( .A(n93), .B(n92), .C(n91), .D(n90), .Y(n94) );
  AOI22XL U245 ( .A(ckcon[0]), .B(n298), .C(dps[0]), .D(n340), .Y(n90) );
  AOI222XL U246 ( .A(ip0[0]), .B(n274), .C(s0rell[0]), .D(n312), .E(ien1[0]), 
        .F(n257), .Y(n93) );
  AOI222XL U247 ( .A(dpc[0]), .B(n261), .C(s0con[0]), .D(n300), .E(s0buf[0]), 
        .F(n297), .Y(n91) );
  AOI221X1 U248 ( .A(tl1[7]), .B(n306), .C(t1_tmod[3]), .D(n305), .E(n304), 
        .Y(n314) );
  AO222XL U249 ( .A(th0[7]), .B(n303), .C(md2[7]), .D(n302), .E(th1[7]), .F(
        n301), .Y(n304) );
  AOI221XL U250 ( .A(s0rell[7]), .B(n312), .C(p2[7]), .D(n311), .E(n310), .Y(
        n313) );
  AO222XL U251 ( .A(sp[7]), .B(n309), .C(dph[7]), .D(n308), .E(dpl[7]), .F(
        n307), .Y(n310) );
  AOI221X1 U252 ( .A(ip0wdts), .B(n274), .C(p2[6]), .D(n311), .E(n273), .Y(
        n275) );
  AO222XL U253 ( .A(dpl[6]), .B(n307), .C(sp[6]), .D(n309), .E(s0rell[6]), .F(
        n312), .Y(n273) );
  AOI222XL U254 ( .A(arcon[0]), .B(n331), .C(b[0]), .D(n332), .E(srstflag), 
        .F(n81), .Y(n84) );
  INVXL U255 ( .A(n80), .Y(n81) );
  AOI222XL U256 ( .A(md3[0]), .B(n289), .C(md4[0]), .D(n291), .E(md5[0]), .F(
        n292), .Y(n83) );
  AOI222XL U257 ( .A(md1[3]), .B(n290), .C(md5[3]), .D(n292), .E(md3[3]), .F(
        n289), .Y(n218) );
  AOI222XL U258 ( .A(md1[1]), .B(n290), .C(md5[1]), .D(n292), .E(md3[1]), .F(
        n289), .Y(n105) );
  AOI222XL U259 ( .A(dph[0]), .B(n308), .C(wdtrel[0]), .D(n293), .E(idle), .F(
        n294), .Y(n87) );
  AOI222XL U260 ( .A(dph[5]), .B(n308), .C(wdtrel[5]), .D(n293), .E(isr_tm), 
        .F(n294), .Y(n263) );
  AOI222XL U261 ( .A(dph[4]), .B(n308), .C(wdtrel[4]), .D(n293), .E(pmw), .F(
        n294), .Y(n240) );
  AOI222XL U262 ( .A(port0[3]), .B(n338), .C(ip1[3]), .D(n249), .E(md0[3]), 
        .F(n329), .Y(n220) );
  AOI222XL U263 ( .A(port0[0]), .B(n338), .C(ip1[0]), .D(n249), .E(md0[0]), 
        .F(n329), .Y(n85) );
  AOI222XL U264 ( .A(port0[1]), .B(n338), .C(ip1[1]), .D(n249), .E(md0[1]), 
        .F(n329), .Y(n107) );
  AOI222XL U265 ( .A(tl1[0]), .B(n306), .C(th0[0]), .D(n303), .E(th1[0]), .F(
        n301), .Y(n89) );
  AOI222XL U266 ( .A(tl1[5]), .B(n306), .C(th0[5]), .D(n303), .E(th1[5]), .F(
        n301), .Y(n265) );
  AOI222XL U267 ( .A(tl1[4]), .B(n306), .C(th0[4]), .D(n303), .E(th1[4]), .F(
        n301), .Y(n242) );
  AOI222XL U268 ( .A(it0), .B(n296), .C(t0_tmod[0]), .D(n305), .E(tl0[0]), .F(
        n295), .Y(n88) );
  AOI222XL U269 ( .A(t0_tf0), .B(n296), .C(t1_tmod[1]), .D(n305), .E(tl0[5]), 
        .F(n295), .Y(n264) );
  AOI222XL U270 ( .A(t0_tr0), .B(n296), .C(t1_tmod[0]), .D(n305), .E(tl0[4]), 
        .F(n295), .Y(n241) );
  AOI222XL U271 ( .A(md4[1]), .B(n291), .C(b[1]), .D(n332), .E(arcon[1]), .F(
        n331), .Y(n106) );
  AOI222XL U272 ( .A(md4[3]), .B(n291), .C(b[3]), .D(n332), .E(arcon[3]), .F(
        n331), .Y(n219) );
  AOI222XL U273 ( .A(ien2[0]), .B(n259), .C(p2[0]), .D(n311), .E(ien0[0]), .F(
        n299), .Y(n92) );
  AO222XL U274 ( .A(s0con[4]), .B(n300), .C(ien2[4]), .D(n259), .E(s0buf[4]), 
        .F(n297), .Y(n238) );
  AO222XL U275 ( .A(s0con[5]), .B(n300), .C(ien2[5]), .D(n259), .E(s0buf[5]), 
        .F(n297), .Y(n260) );
  AO222XL U276 ( .A(ip0[1]), .B(n274), .C(ien1[1]), .D(n257), .E(p2[1]), .F(
        n311), .Y(n101) );
  AO222XL U277 ( .A(ip0[3]), .B(n274), .C(ien1[3]), .D(n257), .E(p2[3]), .F(
        n311), .Y(n214) );
  AO222XL U278 ( .A(md0[5]), .B(n329), .C(ip1[5]), .D(n249), .E(port0[5]), .F(
        n338), .Y(n250) );
  AOI221XL U279 ( .A(dpl[3]), .B(n307), .C(s0rell[3]), .D(n312), .E(n213), .Y(
        n228) );
  AO222XL U280 ( .A(dph[3]), .B(n308), .C(p2sel), .D(n294), .E(sp[3]), .F(n309), .Y(n213) );
  AOI221XL U281 ( .A(dpl[1]), .B(n307), .C(s0rell[1]), .D(n312), .E(n100), .Y(
        n115) );
  AO222XL U282 ( .A(dph[1]), .B(n308), .C(stop), .D(n294), .E(sp[1]), .F(n309), 
        .Y(n100) );
  AO222XL U283 ( .A(i2cadr_o[0]), .B(n323), .C(i2cdat_o[0]), .D(n321), .E(p), 
        .F(n339), .Y(n79) );
  OA21XL U284 ( .B(t1_tr1), .C(t0_tr1), .A(n296), .Y(n279) );
  AOI22XL U285 ( .A(md1[0]), .B(n290), .C(md2[0]), .D(n302), .Y(n82) );
  AOI22XL U286 ( .A(md2[3]), .B(n302), .C(th0[3]), .D(n303), .Y(n217) );
  AOI22XL U287 ( .A(md2[1]), .B(n302), .C(th0[1]), .D(n303), .Y(n104) );
  NOR21XL U288 ( .B(arcon[2]), .A(n171), .Y(n172) );
  NOR21XL U289 ( .B(th0[2]), .A(n159), .Y(n183) );
  NOR21XL U290 ( .B(md2[2]), .A(n160), .Y(n182) );
  NOR21XL U291 ( .B(md4[2]), .A(n170), .Y(n175) );
  NOR21XL U292 ( .B(dpc[2]), .A(n120), .Y(n121) );
  NOR21XL U293 ( .B(ip0[2]), .A(n128), .Y(n137) );
  NOR21XL U294 ( .B(s0buf[2]), .A(n118), .Y(n127) );
  NOR21XL U295 ( .B(ien2[2]), .A(n129), .Y(n136) );
  NOR32XL U296 ( .B(n190), .C(n189), .A(n188), .Y(n208) );
  NOR21XL U297 ( .B(tl1[2]), .A(n187), .Y(n188) );
  NAND21XL U298 ( .B(n186), .A(t0_tmod[2]), .Y(n189) );
  NAND21XL U299 ( .B(n346), .A(th1[2]), .Y(n190) );
  NAND8XL U300 ( .A(n206), .B(n205), .C(n204), .D(n203), .E(n202), .F(n201), 
        .G(n200), .H(n199), .Y(n207) );
  NAND21XL U301 ( .B(n193), .A(dph[2]), .Y(n204) );
  NAND21XL U302 ( .B(n195), .A(dpl[2]), .Y(n202) );
  NAND21XL U303 ( .B(n192), .A(sp[2]), .Y(n205) );
  AO2222XL U304 ( .A(n296), .B(tf1_gate), .C(tl0[7]), .D(n295), .E(smod), .F(
        n294), .G(wdtrel[7]), .H(n293), .Y(n316) );
  AO22XL U305 ( .A(i2cdat_o[2]), .B(n321), .C(ov), .D(n339), .Y(n141) );
  NAND21XL U306 ( .B(n133), .A(ien0[2]), .Y(n134) );
  NAND21XL U307 ( .B(n123), .A(ckcon[2]), .Y(n124) );
  NAND21X1 U308 ( .B(n154), .A(n153), .Y(n155) );
  NOR21XL U309 ( .B(i2ccon_o[2]), .A(n148), .Y(n154) );
  AOI21BBXL U310 ( .B(n152), .C(n151), .A(n150), .Y(n153) );
  NOR21XL U311 ( .B(i2csta_o[2]), .A(n149), .Y(n150) );
  NAND21XL U312 ( .B(n191), .A(gf0), .Y(n206) );
  NAND21XL U313 ( .B(n138), .A(i2cadr_o[2]), .Y(n144) );
  NAND21XL U314 ( .B(n147), .A(s0relh[2]), .Y(n156) );
  NAND21XL U315 ( .B(n140), .A(iex3), .Y(n142) );
  NAND21XL U316 ( .B(n196), .A(tl0[2]), .Y(n201) );
  AND3X1 U317 ( .A(n166), .B(n165), .C(n164), .Y(n181) );
  NAND21XL U318 ( .B(n163), .A(md1[2]), .Y(n164) );
  NAND21XL U319 ( .B(n161), .A(md5[2]), .Y(n166) );
  NAND21XL U320 ( .B(n197), .A(it1), .Y(n200) );
  AOI22XL U321 ( .A(sp[0]), .B(n309), .C(dpl[0]), .D(n307), .Y(n86) );
  AOI22XL U322 ( .A(sp[5]), .B(n309), .C(dpl[5]), .D(n307), .Y(n262) );
  AOI22XL U323 ( .A(sp[4]), .B(n309), .C(dpl[4]), .D(n307), .Y(n239) );
  INVX1 U324 ( .A(acc[2]), .Y(n151) );
  OR2X1 U325 ( .A(t1_tf1), .B(t0_tf1), .Y(tf1_gate) );
  OR2X1 U326 ( .A(s0con[1]), .B(s0con[0]), .Y(riti0_gate) );
  NAND21XL U327 ( .B(n139), .A(t2con[2]), .Y(n143) );
  BUFX3 U328 ( .A(iex2), .Y(iex2_gate) );
  BUFX3 U329 ( .A(iex7), .Y(iex7_gate) );
  BUFX3 U330 ( .A(iex8), .Y(int_vect_8b) );
  BUFX3 U331 ( .A(iex9), .Y(int_vect_93) );
  BUFX3 U332 ( .A(iex10), .Y(int_vect_9b) );
  BUFX3 U333 ( .A(iex11), .Y(int_vect_a3) );
  INVXL U334 ( .A(sfraddr[6]), .Y(n33) );
  INVX1 U335 ( .A(sfraddr[0]), .Y(n26) );
  INVX1 U336 ( .A(n69), .Y(n37) );
  NAND21X1 U337 ( .B(n162), .A(md3[2]), .Y(n165) );
  AND4X2 U338 ( .A(n327), .B(n326), .C(n325), .D(n324), .Y(n334) );
  NOR5X1 U339 ( .A(n309), .B(n308), .C(n307), .D(n257), .E(n312), .Y(n50) );
  AND4X1 U340 ( .A(n256), .B(n255), .C(n254), .D(n253), .Y(n269) );
  NAND21XL U341 ( .B(n194), .A(s0rell[2]), .Y(n203) );
  AOI222XL U342 ( .A(s0relh[7]), .B(n318), .C(port0ff[7]), .D(n341), .E(
        sfrdatai[7]), .F(n317), .Y(n327) );
  AOI222XL U343 ( .A(s0relh[0]), .B(n318), .C(port0ff[0]), .D(n341), .E(
        sfrdatai[0]), .F(n317), .Y(n99) );
  NAND21XL U344 ( .B(n146), .A(sfrdatai[2]), .Y(n157) );
  INVX3 U345 ( .A(n132), .Y(n257) );
  NAND21X2 U346 ( .B(n71), .A(n54), .Y(n132) );
  NAND5X2 U347 ( .A(n345), .B(n347), .C(n77), .D(n343), .E(n342), .Y(n146) );
  NAND6XL U348 ( .A(n347), .B(n346), .C(n345), .D(n344), .E(n343), .F(n342), 
        .Y(ext_sfr_sel) );
  NAND32X1 U349 ( .B(n32), .C(n53), .A(n56), .Y(n47) );
  NAND5XL U350 ( .A(n56), .B(sfraddr[5]), .C(n32), .D(n30), .E(n29), .Y(n130)
         );
  NOR5X1 U351 ( .A(n305), .B(n306), .C(n295), .D(n294), .E(n296), .Y(n72) );
  NAND5XL U352 ( .A(n160), .B(n159), .C(n163), .D(n170), .E(n162), .Y(n73) );
  NAND43X1 U353 ( .B(n75), .C(n74), .D(n73), .A(n72), .Y(n76) );
  AND4X1 U354 ( .A(n224), .B(n223), .C(n222), .D(n221), .Y(n225) );
  NAND6X2 U355 ( .A(n117), .B(n116), .C(n115), .D(n114), .E(n113), .F(n112), 
        .Y(sfrdatao[1]) );
  NAND6X2 U356 ( .A(n248), .B(n247), .C(n246), .D(n245), .E(n244), .F(n243), 
        .Y(sfrdatao[4]) );
  AND4X1 U357 ( .A(n111), .B(n110), .C(n109), .D(n108), .Y(n112) );
  AND4X1 U358 ( .A(n236), .B(n235), .C(n234), .D(n233), .Y(n246) );
  NAND42X4 U359 ( .C(n336), .D(n335), .A(n334), .B(n333), .Y(sfrdatao[7]) );
endmodule


module syncneg_a0 ( clk, reset, rsttowdt, rsttosrst, rst, int0, int1, port0i, 
        rxd0i, sdai, int0ff, int1ff, port0ff, t0ff, t1ff, rxd0ff, sdaiff, 
        rsttowdtff, rsttosrstff, rstff, resetff );
  input [7:0] port0i;
  output [7:0] port0ff;
  input clk, reset, rsttowdt, rsttosrst, rst, int0, int1, rxd0i, sdai;
  output int0ff, int1ff, t0ff, t1ff, rxd0ff, sdaiff, rsttowdtff, rsttosrstff,
         rstff, resetff;
  wire   reset_ff1, int0_ff1, int1_ff1, rxd0_ff1, sdai_ff1;
  wire   [7:0] p0_ff1;

  DFFQX1 reset_ff2_reg ( .D(reset_ff1), .C(clk), .Q(resetff) );
  DFFQX1 rsttosrst_ff1_reg ( .D(rsttosrst), .C(clk), .Q(rsttosrstff) );
  DFFQX1 rsttowdt_ff1_reg ( .D(rsttowdt), .C(clk), .Q(rsttowdtff) );
  DFFQX1 int1_ff2_reg ( .D(int1_ff1), .C(clk), .Q(int1ff) );
  DFFQX1 int0_ff2_reg ( .D(int0_ff1), .C(clk), .Q(int0ff) );
  DFFQX1 rxd0_ff2_reg ( .D(rxd0_ff1), .C(clk), .Q(rxd0ff) );
  DFFQX1 sdai_ff2_reg ( .D(sdai_ff1), .C(clk), .Q(sdaiff) );
  DFFQX1 p0_ff2_reg_7_ ( .D(p0_ff1[7]), .C(clk), .Q(port0ff[7]) );
  DFFQX1 p0_ff2_reg_5_ ( .D(p0_ff1[5]), .C(clk), .Q(port0ff[5]) );
  DFFQX1 p0_ff2_reg_3_ ( .D(p0_ff1[3]), .C(clk), .Q(port0ff[3]) );
  DFFQX1 p0_ff2_reg_1_ ( .D(p0_ff1[1]), .C(clk), .Q(port0ff[1]) );
  DFFQX1 p0_ff2_reg_0_ ( .D(p0_ff1[0]), .C(clk), .Q(port0ff[0]) );
  DFFQX1 p0_ff2_reg_6_ ( .D(p0_ff1[6]), .C(clk), .Q(port0ff[6]) );
  DFFQX1 p0_ff2_reg_2_ ( .D(p0_ff1[2]), .C(clk), .Q(port0ff[2]) );
  DFFQX1 p0_ff2_reg_4_ ( .D(p0_ff1[4]), .C(clk), .Q(port0ff[4]) );
  DFFQX1 rst_ff1_reg ( .D(rst), .C(clk), .Q(rstff) );
  DFFQX1 int0_ff1_reg ( .D(int0), .C(clk), .Q(int0_ff1) );
  DFFQX1 int1_ff1_reg ( .D(int1), .C(clk), .Q(int1_ff1) );
  DFFQX1 p0_ff1_reg_6_ ( .D(port0i[6]), .C(clk), .Q(p0_ff1[6]) );
  DFFQX1 p0_ff1_reg_5_ ( .D(port0i[5]), .C(clk), .Q(p0_ff1[5]) );
  DFFQX1 p0_ff1_reg_4_ ( .D(port0i[4]), .C(clk), .Q(p0_ff1[4]) );
  DFFQX1 p0_ff1_reg_2_ ( .D(port0i[2]), .C(clk), .Q(p0_ff1[2]) );
  DFFQX1 p0_ff1_reg_1_ ( .D(port0i[1]), .C(clk), .Q(p0_ff1[1]) );
  DFFQX1 p0_ff1_reg_0_ ( .D(port0i[0]), .C(clk), .Q(p0_ff1[0]) );
  DFFQX1 rxd0_ff1_reg ( .D(rxd0i), .C(clk), .Q(rxd0_ff1) );
  DFFQX1 p0_ff1_reg_7_ ( .D(port0i[7]), .C(clk), .Q(p0_ff1[7]) );
  DFFQX1 p0_ff1_reg_3_ ( .D(port0i[3]), .C(clk), .Q(p0_ff1[3]) );
  DFFQX1 sdai_ff1_reg ( .D(sdai), .C(clk), .Q(sdai_ff1) );
  DFFQX1 reset_ff1_reg ( .D(reset), .C(clk), .Q(reset_ff1) );
  INVX1 U3 ( .A(1'b1), .Y(t1ff) );
  INVX1 U5 ( .A(1'b1), .Y(t0ff) );
endmodule


module mcu51_cpu_a0 ( clkcpu, rst, mempsack, memack, memdatai, memaddr, 
        mempsrd, mempswr, memrd, memwr, memaddr_comb, mempsrd_comb, 
        mempswr_comb, memrd_comb, memwr_comb, cpu_hold, cpu_resume, irq, 
        intvect, intcall, retiinstr, newinstr, rmwinstr, waitstaten, ramdatai, 
        sfrdatai, ramsfraddr, ramdatao, ramoe, ramwe, sfroe, sfrwe, sfroe_r, 
        sfrwe_r, sfroe_comb_s, sfrwe_comb_s, pc_o, pc_ini, cs_run, instr, 
        codefetch_s, sfrack, ramsfraddr_comb, ramdatao_comb, ramoe_comb, 
        ramwe_comb, ckcon, pmw, p2sel, gf0, stop, idle, acc, b, rs, c, ac, ov, 
        p, f0, f1, dph, dpl, dps, dpc, p2, sp );
  input [7:0] memdatai;
  output [15:0] memaddr;
  output [15:0] memaddr_comb;
  input [4:0] intvect;
  input [7:0] ramdatai;
  input [7:0] sfrdatai;
  output [7:0] ramsfraddr;
  output [7:0] ramdatao;
  output [15:0] pc_o;
  input [15:0] pc_ini;
  output [7:0] instr;
  output [7:0] ramsfraddr_comb;
  output [7:0] ramdatao_comb;
  output [7:0] ckcon;
  output [7:0] acc;
  output [7:0] b;
  output [1:0] rs;
  output [7:0] dph;
  output [7:0] dpl;
  output [3:0] dps;
  output [5:0] dpc;
  output [7:0] p2;
  output [7:0] sp;
  input clkcpu, rst, mempsack, memack, cpu_hold, cpu_resume, irq, sfrack;
  output mempsrd, mempswr, memrd, memwr, mempsrd_comb, mempswr_comb,
         memrd_comb, memwr_comb, intcall, retiinstr, newinstr, rmwinstr,
         waitstaten, ramoe, ramwe, sfroe, sfrwe, sfroe_r, sfrwe_r,
         sfroe_comb_s, sfrwe_comb_s, cs_run, codefetch_s, ramoe_comb,
         ramwe_comb, pmw, p2sel, gf0, stop, idle, c, ac, ov, p, f0, f1;
  wire   N343, N344, N345, N346, N347, N348, N350, N352, N353, N354, n2184,
         n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194,
         finishmul, finishdiv, N370, N371, N372, N480, N481, N482, N483, N484,
         N485, N486, N487, N488, N489, N490, N491, N492, N493, N494, N495,
         d_hold, idle_r, cpu_resume_fff, stop_r, ramsfrwe, N512, N515, N520,
         pdmode, interrupt, N582, N583, N584, N585, N588, N589, N590,
         phase0_ff, newinstrlock, N670, N671, N672, N673, N674, N675, N676,
         N677, N679, N680, N681, N682, N683, N684, N685, N689, N690, N1761,
         N1763, N1764, N1765, N1766, N1767, N1768, accactv, N10562, N10563,
         N10564, N10565, N10566, N10567, N10568, N10569, N10570, N10571,
         N10572, N10573, N10574, N10575, N10576, N10577, N10578, N10579,
         N10580, N10581, N10582, N10583, N10584, N10585, N10586, N10587,
         N10588, N10589, N11478, N11479, N11480, N11481, N11482, N11483,
         N11484, N11485, N11486, N11487, N11488, N11489, N11491, N11492,
         N11493, N11494, N11498, N11499, N11500, N11501, N11502, N11503,
         N11504, N11505, N11522, N11523, N11524, N11525, N11526, N11527,
         N11528, N11541, N11542, N11543, N11544, N11545, N11546, N11547,
         N11549, N11555, N11560, N11584, N11780, N11781, N11782, N11783,
         N11784, N11785, N11786, N11787, N11788, N11789, N11790, N11791,
         N11792, N11793, N11796, N11797, N11798, N11799, N11800, N11801,
         N11802, N11803, N11804, N11805, N11806, N11807, N11808, N11809,
         N11810, N11814, N11815, N11816, N11817, N11818, N11819, N11820,
         N11821, N11822, N11823, N11824, N11825, N11826, N11827, N11835,
         N11836, N11837, N11838, N11839, N11840, N11841, N11842, N11845,
         N11846, N11847, N11848, N11849, N11850, N11851, N11852, N12469,
         N12470, N12471, N12472, N12473, N12474, N12475, N12476, N12477,
         N12478, N12479, N12480, N12481, N12482, N12483, N12484, N12485,
         N12486, N12487, N12488, N12489, N12490, N12491, N12492, N12493,
         N12494, N12495, N12496, N12497, N12498, N12499, N12500, N12501,
         N12502, N12503, N12504, N12505, N12506, N12507, N12508, N12509,
         N12510, N12511, N12512, N12513, N12514, N12515, N12516, N12517,
         N12518, N12519, N12520, N12521, N12522, N12523, N12524, N12525,
         N12526, N12527, N12528, N12529, N12530, N12531, N12532, N12533,
         N12534, N12535, N12536, N12537, N12538, N12539, N12540, N12541,
         N12542, N12543, N12544, N12545, N12546, N12547, N12548, N12549,
         N12550, N12551, N12552, N12553, N12554, N12555, N12556, N12557,
         N12558, N12559, N12560, N12561, N12562, N12563, N12564, N12566,
         N12567, N12568, N12569, N12570, N12571, N12572, N12573, N12575,
         N12576, N12577, N12578, N12579, N12580, N12581, N12582, N12584,
         N12585, N12586, N12587, N12588, N12589, N12590, N12591, N12593,
         N12594, N12595, N12596, N12597, N12598, N12599, N12600, N12602,
         N12603, N12604, N12605, N12606, N12607, N12608, N12609, N12611,
         N12612, N12613, N12614, N12615, N12616, N12617, N12618, N12620,
         N12621, N12622, N12623, N12624, N12625, N12626, N12627, N12629,
         N12630, N12631, N12632, N12633, N12634, N12635, N12636, N12637,
         N12644, N12651, N12658, N12665, N12672, N12679, N12686, N12690,
         N12691, N12692, N12693, N12694, N12695, N12697, N12698, N12699,
         N12700, N12701, N12702, N12703, N12704, N12705, N12706, N12709,
         N12710, N12711, N12714, N12715, N12716, N12717, N12718, N12719,
         N12720, N12721, N12722, N12723, N12724, N12725, N12726, N12727,
         N12728, N12729, N12730, N12769, N12770, N12771, N12772, N12773,
         N12774, N12775, N12776, N12801, N12802, N12803, N12804, N12805,
         N12806, N12807, N12808, N12810, N12811, N12812, N12813, N12814,
         N12815, N12816, N12817, N12824, N12825, N12826, N12827, N12828,
         N12829, N12830, N12831, N12841, N12842, N12843, N12844, N12845,
         N12846, N12847, N12848, N12849, N12850, N12851, N12852, N12853,
         N12854, N12855, N12856, N12905, israccess, N12912, N12965, N12966,
         N12967, N12968, N12969, N12970, N12971, N12972, N12974, N12975,
         N12976, N12977, N13014, N13023, N13032, N13041, N13050, N13059,
         N13068, N13077, N13086, N13095, N13104, N13113, N13122, N13131,
         N13140, N13149, N13158, N13167, N13176, N13185, N13194, N13203,
         N13212, N13221, N13230, N13239, N13248, N13257, N13266, N13275,
         N13284, N13293, multemp1_0_, N13324, N13325, N13326, N13327, N13328,
         N13329, N13330, N13331, N13332, N13336, N13337, N13338, N13339,
         N13340, N13341, N13342, N13343, divtemp1_0_, N13345, N13346, N13347,
         N13348, N13349, N13350, N13351, N13352, N13353, N13366, N13367,
         N13368, N13369, N13370, N13371, N13372, N13373, cpu_resume_ff1,
         N13379, N13380, net12400, net12406, net12411, net12416, net12421,
         net12426, net12431, net12436, net12441, net12446, net12451, net12456,
         net12461, net12466, net12471, net12476, net12481, net12486, net12491,
         net12496, net12501, net12506, net12511, net12516, net12521, net12526,
         net12531, net12536, net12541, net12546, net12551, net12556, net12561,
         net12566, net12571, net12576, net12581, net12586, net12591, net12596,
         net12601, net12606, net12611, net12616, net12621, net12626, net12631,
         net12636, net12641, net12646, net12651, net12656, net12661, net12666,
         net12671, n658, n661, n662, n667, n670, n671, n672, n673, n678, n680,
         n681, n683, n684, n685, n686, n687, n688, n693, n695, n696, n716,
         n717, n719, n720, n721, n722, n723, n725, n726, n727, n730, n733,
         n734, n736, n737, n742, n743, n744, n745, n747, n748, n749, n750,
         n751, n757, n763, n775, n780, n785, n790, n795, n801, n807, n812,
         n817, n836, n841, n842, n847, n848, n853, n854, n860, n865, n866,
         n871, n872, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n926, n929, n930, n931, n932, n933, n940, n949,
         n960, n964, n967, n968, n969, n970, n972, n977, n978, n998, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1023, n1024, n1025, n1029, n1030, n1031,
         n1032, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1048, n1051, n1053, n1054, n1055, n1056,
         n1057, n1061, n1062, n1063, n1066, n1067, n1068, n1069, n1070, n1071,
         n1072, n1073, n1076, n1077, n1080, n1081, n1084, n1085, n1088, n1089,
         n1090, n1092, n1093, n1094, n1096, n1097, n1098, n1100, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1150, n1151, n1152, n1153, n1154, n1155,
         n1156, n1157, n1158, n1159, n1162, n1163, n1164, n1165, n1166, n1167,
         n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
         n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
         n1188, n1189, n1190, n1191, n1192, n1194, n1195, n1196, n1199, n1200,
         n1201, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
         n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
         n1222, n1223, n1224, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
         n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
         n1266, n1267, n1268, n1269, n1270, n1271, n1275, n1276, n1277, n1278,
         n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
         n1289, n1305, n1306, n1307, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1323, n1324, n1325,
         n1326, n1327, n1328, n1329, n1331, n1332, n1333, n1335, n1336, n1337,
         n1338, n1339, n1340, n1341, n1342, n1345, n1346, n1347, n1348, n1349,
         n1355, n1356, n1357, n1358, n1360, n1363, n1364, n1365, n1366, n1369,
         n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
         n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1391, n1392,
         n1393, n1394, n1395, n1397, n1398, n1400, n1403, n1405, n1406, n1407,
         n1408, n1409, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
         n1430, n1431, n1435, n1436, n1437, n1445, n1446, n1447, n1448, n1449,
         n1456, n1457, n1458, n1462, n1463, n1464, n1465, n1466, n1467, n1468,
         n1470, n1471, n1472, n1473, n1480, n1482, n1486, n1487, n1488, n1489,
         n1490, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1513,
         n1514, n1516, n1517, n1518, n1520, n1531, n1532, n1549, n1550, n1573,
         n1575, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1585, n1586,
         n1589, n1590, n1591, n1593, n1594, n1597, n1598, n1599, n1600, n1601,
         n1602, n1605, n1608, n1609, n1611, n1614, n1618, n1619, n1620, n1622,
         n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1633, n1635,
         n1636, n1637, n1638, n1639, n1640, n1647, n1648, n1649, n1650, n1651,
         n1652, n1653, n1654, n1657, n1658, n1660, n1662, n1667, n1668, n1669,
         n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679,
         n1680, n1681, n1682, n1683, n1685, n1686, n1687, n1688, n1689, n1691,
         n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701,
         n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1723,
         n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733,
         n1734, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
         n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
         n1755, n1756, n1758, n1760, n1761, n1762, n1764, n1765, n1766, n1767,
         n1768, n1769, n1770, n1771, n1772, n1774, n1775, n1776, n1777, n1778,
         n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788,
         n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798,
         n1799, n1800, n1801, n1802, n1803, n1805, n1806, n1807, n1809, n1810,
         n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820,
         n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830,
         n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, multemp1_8_, multemp1_7_, multemp1_6_, multemp1_5_,
         multemp1_4_, multemp1_3_, multemp1_2_, multemp1_1_, N14351, N14350,
         N14349, N14348, N14347, N14346, N14345, N14344, N14343, N14342,
         N14341, N14340, N14339, N14338, N14337, N14336, add_5526_carry_2_,
         add_5526_carry_3_, add_5526_carry_4_, add_5526_carry_5_,
         add_5526_carry_6_, add_5526_carry_7_, add_5280_3_carry_2_,
         add_5280_3_carry_3_, add_5280_3_carry_4_, add_5280_3_carry_5_,
         add_5280_3_carry_6_, add_5280_3_carry_7_, add_5280_3_carry_8_,
         add_5280_3_carry_9_, add_5280_3_carry_10_, add_5280_3_carry_11_,
         add_5280_3_carry_12_, add_5280_3_carry_13_, add_5280_3_carry_14_,
         add_5280_3_carry_15_, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n19, n21, n22, n23, n25, n27, n29, n31, n33, n35, n37,
         n39, n41, n43, n45, n47, n49, n50, n53, n56, n57, n58, n60, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n123, n124, n125, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n440, n441,
         n442, n444, n445, n446, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n659, n660, n663, n664, n665, n666,
         n668, n669, n674, n675, n676, n677, n679, n682, n689, n690, n691,
         n692, n694, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n718,
         n724, n728, n729, n731, n732, n735, n738, n739, n740, n741, n746,
         n752, n753, n754, n755, n756, n758, n759, n760, n761, n762, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n776,
         n777, n778, n779, n781, n782, n783, n784, n786, n787, n788, n789,
         n791, n792, n793, n794, n796, n797, n798, n799, n800, n802, n803,
         n804, n805, n806, n808, n809, n810, n811, n813, n814, n815, n816,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n837, n838, n839, n840,
         n843, n844, n845, n846, n849, n850, n851, n852, n855, n856, n857,
         n858, n859, n861, n862, n863, n864, n867, n868, n869, n870, n873,
         n874, n875, n876, n877, n878, n879, n925, n927, n928, n934, n935,
         n936, n937, n938, n939, n941, n942, n943, n944, n945, n946, n947,
         n948, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n961, n962, n963, n965, n966, n971, n973, n974, n975, n976, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n999, n1008, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1026, n1027, n1028, n1033, n1047,
         n1049, n1050, n1052, n1058, n1059, n1060, n1064, n1065, n1074, n1075,
         n1078, n1079, n1082, n1083, n1086, n1087, n1091, n1095, n1099, n1101,
         n1131, n1149, n1160, n1161, n1193, n1197, n1198, n1202, n1225, n1233,
         n1234, n1248, n1272, n1273, n1274, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1308, n1322, n1330, n1334, n1343, n1344, n1350, n1351, n1352, n1353,
         n1354, n1359, n1361, n1362, n1367, n1368, n1388, n1389, n1390, n1396,
         n1399, n1401, n1402, n1404, n1410, n1411, n1412, n1413, n1414, n1415,
         n1416, n1417, n1418, n1419, n1420, n1421, n1432, n1433, n1434, n1438,
         n1439, n1440, n1441, n1442, n1443, n1444, n1450, n1451, n1452, n1453,
         n1454, n1455, n1459, n1460, n1461, n1469, n1474, n1475, n1476, n1477,
         n1478, n1479, n1481, n1483, n1484, n1485, n1491, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1515, n1519, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528,
         n1529, n1530, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540,
         n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1574, n1576, n1584, n1587, n1588, n1592, n1595, n1596, n1603, n1604,
         n1606, n1607, n1610, n1612, n1613, n1615, n1616, n1617, n1621, n1623,
         n1632, n1634, n1641, n1642, n1643, n1644, n1645, n1646, n1655, n1656,
         n1659, n1661, n1663, n1664, n1665, n1666, n1684, n1690, n1710, n1722,
         n1735, n1757, n1759, n1763, n1773, n1804, n1808, n1840, n1841, n1885,
         n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895,
         n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905,
         n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915,
         n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925,
         n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935,
         n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945,
         n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955,
         n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965,
         n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975,
         n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985,
         n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995,
         n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005,
         n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015,
         n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025,
         n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035,
         n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045,
         n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055,
         n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065,
         n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075,
         n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085,
         n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095,
         n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105,
         n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115,
         n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125,
         n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135,
         n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145,
         n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155,
         n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165,
         n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2177, n2178,
         n2179, n2180, n2181, n2182, n2183, SYNOPSYS_UNCONNECTED_1;
  wire   [2:0] state;
  wire   [5:0] phase;
  wire   [15:0] alu_out;
  wire   [15:0] pc_i;
  wire   [7:0] temp;
  wire   [7:4] incdec_out;
  wire   [18:0] dec_accop;
  wire   [7:0] dec_cop;
  wire   [6:2] adder_out;
  wire   [9:1] multemp2;
  wire   [7:0] temp2_comb;
  wire   [7:0] dph_current;
  wire   [7:0] dpl_current;
  wire   [15:0] dptr_inc;
  wire   [63:0] dpl_reg;
  wire   [63:0] dph_reg;
  wire   [47:0] dpc_tab;
  wire   [2:0] waitcnt;
  wire   [255:0] rn_reg;
  wire   [6:0] rn;
  wire   [7:0] multempreg;
  wire   [6:0] divtempreg;
  wire   [15:3] add_5280_4_carry;
  wire   [15:3] add_5280_2_carry;
  wire   [7:3] add_1469_carry;
  wire   [3:2] add_1_root_add_5140_2_carry;

  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_0 clk_gate_finishmul_reg ( .CLK(clkcpu), 
        .EN(N370), .ENCLK(net12400), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_54 clk_gate_instr_reg ( .CLK(clkcpu), .EN(
        N685), .ENCLK(net12406), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_53 clk_gate_bitno_reg ( .CLK(clkcpu), .EN(
        N11491), .ENCLK(net12411), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_52 clk_gate_dph_reg_reg_7_ ( .CLK(clkcpu), 
        .EN(N12556), .ENCLK(net12416), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_51 clk_gate_dph_reg_reg_6_ ( .CLK(clkcpu), 
        .EN(N12547), .ENCLK(net12421), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_50 clk_gate_dph_reg_reg_5_ ( .CLK(clkcpu), 
        .EN(N12538), .ENCLK(net12426), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_49 clk_gate_dph_reg_reg_4_ ( .CLK(clkcpu), 
        .EN(N12529), .ENCLK(net12431), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_48 clk_gate_dph_reg_reg_3_ ( .CLK(clkcpu), 
        .EN(N12520), .ENCLK(net12436), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_47 clk_gate_dph_reg_reg_2_ ( .CLK(clkcpu), 
        .EN(N12511), .ENCLK(net12441), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_46 clk_gate_dph_reg_reg_1_ ( .CLK(clkcpu), 
        .EN(N12502), .ENCLK(net12446), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_45 clk_gate_dph_reg_reg_0_ ( .CLK(clkcpu), 
        .EN(N12493), .ENCLK(net12451), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_44 clk_gate_dpc_tab_reg_7_ ( .CLK(clkcpu), 
        .EN(N12686), .ENCLK(net12456), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_43 clk_gate_dpc_tab_reg_6_ ( .CLK(clkcpu), 
        .EN(N12679), .ENCLK(net12461), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_42 clk_gate_dpc_tab_reg_5_ ( .CLK(clkcpu), 
        .EN(N12672), .ENCLK(net12466), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_41 clk_gate_dpc_tab_reg_4_ ( .CLK(clkcpu), 
        .EN(N12665), .ENCLK(net12471), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_40 clk_gate_dpc_tab_reg_3_ ( .CLK(clkcpu), 
        .EN(N12658), .ENCLK(net12476), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_39 clk_gate_dpc_tab_reg_2_ ( .CLK(clkcpu), 
        .EN(N12651), .ENCLK(net12481), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_38 clk_gate_dpc_tab_reg_1_ ( .CLK(clkcpu), 
        .EN(N12644), .ENCLK(net12486), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_37 clk_gate_dpc_tab_reg_0_ ( .CLK(clkcpu), 
        .EN(N12637), .ENCLK(net12491), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_36 clk_gate_temp_reg ( .CLK(clkcpu), .EN(
        N12722), .ENCLK(net12496), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_35 clk_gate_waitcnt_reg ( .CLK(clkcpu), 
        .EN(N12977), .ENCLK(net12501), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_34 clk_gate_rn_reg_reg_0_ ( .CLK(clkcpu), 
        .EN(N13293), .ENCLK(net12506), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_33 clk_gate_rn_reg_reg_1_ ( .CLK(clkcpu), 
        .EN(N13284), .ENCLK(net12511), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_32 clk_gate_rn_reg_reg_2_ ( .CLK(clkcpu), 
        .EN(N13275), .ENCLK(net12516), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_31 clk_gate_rn_reg_reg_3_ ( .CLK(clkcpu), 
        .EN(N13266), .ENCLK(net12521), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_30 clk_gate_rn_reg_reg_4_ ( .CLK(clkcpu), 
        .EN(N13257), .ENCLK(net12526), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_29 clk_gate_rn_reg_reg_5_ ( .CLK(clkcpu), 
        .EN(N13248), .ENCLK(net12531), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_28 clk_gate_rn_reg_reg_6_ ( .CLK(clkcpu), 
        .EN(N13239), .ENCLK(net12536), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_27 clk_gate_rn_reg_reg_7_ ( .CLK(clkcpu), 
        .EN(N13230), .ENCLK(net12541), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_26 clk_gate_rn_reg_reg_8_ ( .CLK(clkcpu), 
        .EN(N13221), .ENCLK(net12546), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_25 clk_gate_rn_reg_reg_9_ ( .CLK(clkcpu), 
        .EN(N13212), .ENCLK(net12551), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_24 clk_gate_rn_reg_reg_10_ ( .CLK(clkcpu), 
        .EN(N13203), .ENCLK(net12556), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_23 clk_gate_rn_reg_reg_11_ ( .CLK(clkcpu), 
        .EN(N13194), .ENCLK(net12561), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_22 clk_gate_rn_reg_reg_12_ ( .CLK(clkcpu), 
        .EN(N13185), .ENCLK(net12566), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_21 clk_gate_rn_reg_reg_13_ ( .CLK(clkcpu), 
        .EN(N13176), .ENCLK(net12571), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_20 clk_gate_rn_reg_reg_14_ ( .CLK(clkcpu), 
        .EN(N13167), .ENCLK(net12576), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_19 clk_gate_rn_reg_reg_15_ ( .CLK(clkcpu), 
        .EN(N13158), .ENCLK(net12581), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_18 clk_gate_rn_reg_reg_16_ ( .CLK(clkcpu), 
        .EN(N13149), .ENCLK(net12586), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_17 clk_gate_rn_reg_reg_17_ ( .CLK(clkcpu), 
        .EN(N13140), .ENCLK(net12591), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_16 clk_gate_rn_reg_reg_18_ ( .CLK(clkcpu), 
        .EN(N13131), .ENCLK(net12596), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_15 clk_gate_rn_reg_reg_19_ ( .CLK(clkcpu), 
        .EN(N13122), .ENCLK(net12601), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_14 clk_gate_rn_reg_reg_20_ ( .CLK(clkcpu), 
        .EN(N13113), .ENCLK(net12606), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_13 clk_gate_rn_reg_reg_21_ ( .CLK(clkcpu), 
        .EN(N13104), .ENCLK(net12611), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_12 clk_gate_rn_reg_reg_22_ ( .CLK(clkcpu), 
        .EN(N13095), .ENCLK(net12616), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_11 clk_gate_rn_reg_reg_23_ ( .CLK(clkcpu), 
        .EN(N13086), .ENCLK(net12621), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_10 clk_gate_rn_reg_reg_24_ ( .CLK(clkcpu), 
        .EN(N13077), .ENCLK(net12626), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_9 clk_gate_rn_reg_reg_25_ ( .CLK(clkcpu), 
        .EN(N13068), .ENCLK(net12631), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_8 clk_gate_rn_reg_reg_26_ ( .CLK(clkcpu), 
        .EN(N13059), .ENCLK(net12636), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_7 clk_gate_rn_reg_reg_27_ ( .CLK(clkcpu), 
        .EN(N13050), .ENCLK(net12641), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_6 clk_gate_rn_reg_reg_28_ ( .CLK(clkcpu), 
        .EN(N13041), .ENCLK(net12646), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_5 clk_gate_rn_reg_reg_29_ ( .CLK(clkcpu), 
        .EN(N13032), .ENCLK(net12651), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_4 clk_gate_rn_reg_reg_30_ ( .CLK(clkcpu), 
        .EN(N13023), .ENCLK(net12656), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_3 clk_gate_rn_reg_reg_31_ ( .CLK(clkcpu), 
        .EN(N13014), .ENCLK(net12661), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_2 clk_gate_multempreg_reg ( .CLK(clkcpu), 
        .EN(N13324), .ENCLK(net12666), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_1 clk_gate_divtempreg_reg ( .CLK(clkcpu), 
        .EN(N13366), .ENCLK(net12671), .TE(1'b0) );
  mcu51_cpu_a0_DW01_add_0 add_5586 ( .A({n1894, n1894, n1894, n1894, n1894, 
        n1894, n1894, n1894, N12831, N12830, N12829, N12828, N12827, N12826, 
        N12825, N12824}), .B({N12856, N12855, N12854, N12853, N12852, N12851, 
        N12850, N12849, N12848, N12847, N12846, N12845, N12844, N12843, N12842, 
        N12841}), .CI(1'b0), .SUM(alu_out), .CO() );
  mcu51_cpu_a0_DW01_sub_0 sub_5969 ( .A({1'b0, n189, n188, n187, n186, n185, 
        n184, divtemp1_0_, acc[6]}), .B({1'b0, b}), .CI(1'b0), .DIFF({N13353, 
        N13352, N13351, N13350, N13349, N13348, N13347, N13346, N13345}), 
        .CO() );
  mcu51_cpu_a0_DW01_sub_1 sub_5950 ( .A({1'b0, divtempreg, n70}), .B({1'b0, b}), .CI(1'b0), .DIFF({N13343, SYNOPSYS_UNCONNECTED_1, N13342, N13341, N13340, 
        N13339, N13338, N13337, N13336}), .CO() );
  mcu51_cpu_a0_DW01_inc_0 add_5525 ( .A({N12776, N12775, N12774, N12773, 
        N12772, N12771, N12770, N12769}), .SUM({N12808, N12807, N12806, N12805, 
        N12804, N12803, N12802, N12801}) );
  mcu51_cpu_a0_DW01_inc_1 add_5286 ( .A({dph_current, dpl_current}), .SUM(
        dptr_inc) );
  mcu51_cpu_a0_DW01_inc_2 r715 ( .A({pc_o[15:14], n49, pc_o[12:7], 
        memaddr[6:5], pc_o[4:0]}), .SUM(pc_i) );
  mcu51_cpu_a0_DW01_add_8 add_5901_aco ( .A({1'b0, multempreg}), .B({1'b0, 
        N14343, N14342, N14341, N14340, N14339, N14338, N14337, N14336}), .CI(
        1'b0), .SUM({multemp1_8_, multemp1_7_, multemp1_6_, multemp1_5_, 
        multemp1_4_, multemp1_3_, multemp1_2_, multemp1_1_, multemp1_0_}), 
        .CO() );
  mcu51_cpu_a0_DW01_add_7 add_5907_aco ( .A({1'b0, multemp1_8_, multemp1_7_, 
        multemp1_6_, multemp1_5_, multemp1_4_, multemp1_3_, multemp1_2_, 
        multemp1_1_}), .B({1'b0, N14351, N14350, N14349, N14348, N14347, 
        N14346, N14345, N14344}), .CI(1'b0), .SUM(multemp2), .CO() );
  FAD1X1 add_1_root_add_5140_2_U1_2 ( .A(N11524), .B(N11543), .CI(
        add_1_root_add_5140_2_carry[2]), .CO(add_1_root_add_5140_2_carry[3]), 
        .SO(adder_out[2]) );
  FAD1X1 add_1_root_add_5140_2_U1_3 ( .A(N11525), .B(N11544), .CI(
        add_1_root_add_5140_2_carry[3]), .CO(N11555), .SO(adder_out[3]) );
  DFFQX1 cpu_resume_ff1_reg ( .D(N13379), .C(clkcpu), .Q(cpu_resume_ff1) );
  DFFQX1 newinstrlock_reg ( .D(n1878), .C(net12400), .Q(newinstrlock) );
  DFFQX1 phase0_ff_reg ( .D(N689), .C(net12400), .Q(phase0_ff) );
  DFFQX1 finishdiv_reg ( .D(N372), .C(net12400), .Q(finishdiv) );
  DFFQX1 finishmul_reg ( .D(N371), .C(net12400), .Q(finishmul) );
  DFFQX1 multempreg_reg_7_ ( .D(N13332), .C(net12666), .Q(multempreg[7]) );
  DFFQX1 multempreg_reg_6_ ( .D(N13331), .C(net12666), .Q(multempreg[6]) );
  DFFQX1 multempreg_reg_5_ ( .D(N13330), .C(net12666), .Q(multempreg[5]) );
  DFFQX1 pdmode_reg ( .D(n1973), .C(net12400), .Q(pdmode) );
  DFFQX1 multempreg_reg_4_ ( .D(N13329), .C(net12666), .Q(multempreg[4]) );
  DFFQX1 d_hold_reg ( .D(cpu_hold), .C(clkcpu), .Q(d_hold) );
  DFFQX1 cpu_resume_fff_reg ( .D(N13380), .C(clkcpu), .Q(cpu_resume_fff) );
  DFFQX1 multempreg_reg_3_ ( .D(N13328), .C(net12666), .Q(multempreg[3]) );
  DFFQX1 multempreg_reg_2_ ( .D(N13327), .C(net12666), .Q(multempreg[2]) );
  DFFQX1 idle_r_reg ( .D(N512), .C(net12400), .Q(idle_r) );
  DFFQX1 stop_r_reg ( .D(N515), .C(net12400), .Q(stop_r) );
  DFFQX1 ramoe_r_reg ( .D(N11486), .C(net12400), .Q(ramoe) );
  DFFQX1 phase_reg_5_ ( .D(N684), .C(net12400), .Q(phase[5]) );
  DFFQX1 state_reg_1_ ( .D(N589), .C(net12400), .Q(state[1]) );
  DFFQX1 state_reg_2_ ( .D(N590), .C(net12400), .Q(state[2]) );
  DFFQX1 israccess_reg ( .D(N12912), .C(net12400), .Q(israccess) );
  DFFQX1 phase_reg_4_ ( .D(N683), .C(net12400), .Q(phase[4]) );
  DFFQX1 state_reg_0_ ( .D(N588), .C(net12400), .Q(state[0]) );
  DFFQX1 phase_reg_3_ ( .D(N682), .C(net12400), .Q(phase[3]) );
  DFFQX1 dec_cop_reg_0_ ( .D(N10582), .C(net12400), .Q(dec_cop[0]) );
  DFFQX1 f0_reg ( .D(n1882), .C(net12400), .Q(f0) );
  DFFQX1 ov_reg_reg ( .D(N12711), .C(net12400), .Q(ov) );
  DFFQX1 gf0_reg ( .D(n1881), .C(net12400), .Q(gf0) );
  DFFQX1 p2_reg_reg_7_ ( .D(N12492), .C(net12400), .Q(p2[7]) );
  DFFQX1 p2_reg_reg_5_ ( .D(N12490), .C(net12400), .Q(p2[5]) );
  DFFQX1 p2_reg_reg_4_ ( .D(N12489), .C(net12400), .Q(p2[4]) );
  DFFQX1 dpc_tab_reg_3__5_ ( .D(n409), .C(net12476), .Q(dpc_tab[23]) );
  DFFQX1 dpc_tab_reg_3__4_ ( .D(N12691), .C(net12476), .Q(dpc_tab[22]) );
  DFFQX1 dpc_tab_reg_7__5_ ( .D(N12692), .C(net12456), .Q(dpc_tab[47]) );
  DFFQX1 dpc_tab_reg_0__5_ ( .D(n410), .C(net12491), .Q(dpc_tab[5]) );
  DFFQX1 dpc_tab_reg_0__4_ ( .D(n412), .C(net12491), .Q(dpc_tab[4]) );
  DFFQX1 dpc_tab_reg_4__5_ ( .D(N12692), .C(net12471), .Q(dpc_tab[29]) );
  DFFQX1 dpc_tab_reg_1__5_ ( .D(n409), .C(net12486), .Q(dpc_tab[11]) );
  DFFQX1 dpc_tab_reg_2__5_ ( .D(n409), .C(net12481), .Q(dpc_tab[17]) );
  DFFQX1 dpc_tab_reg_2__4_ ( .D(N12691), .C(net12481), .Q(dpc_tab[16]) );
  DFFQX1 dpc_tab_reg_6__5_ ( .D(N12692), .C(net12461), .Q(dpc_tab[41]) );
  DFFQX1 p_reg ( .D(N12905), .C(net12400), .Q(p) );
  DFFQX1 dec_cop_reg_5_ ( .D(N10587), .C(net12400), .Q(dec_cop[5]) );
  DFFQX1 dec_cop_reg_2_ ( .D(N10584), .C(net12400), .Q(dec_cop[2]) );
  DFFQX1 sp_reg_reg_7_ ( .D(N12704), .C(net12400), .Q(sp[7]) );
  DFFQX1 dpl_reg_reg_3__3_ ( .D(N12596), .C(net12436), .Q(dpl_reg[27]) );
  DFFQX1 dpl_reg_reg_0__3_ ( .D(N12569), .C(net12451), .Q(dpl_reg[3]) );
  DFFQX1 dpl_reg_reg_2__3_ ( .D(N12587), .C(net12441), .Q(dpl_reg[19]) );
  DFFQX1 dec_cop_reg_3_ ( .D(N10585), .C(net12400), .Q(dec_cop[3]) );
  DFFQX1 dec_cop_reg_1_ ( .D(N10583), .C(net12400), .Q(dec_cop[1]) );
  DFFQX1 dec_cop_reg_4_ ( .D(N10586), .C(net12400), .Q(dec_cop[4]) );
  DFFQX1 multempreg_reg_1_ ( .D(N13326), .C(net12666), .Q(multempreg[1]) );
  DFFQX1 p2sel_s_reg ( .D(N520), .C(net12400), .Q(p2sel) );
  DFFQX1 p2_reg_reg_1_ ( .D(N12486), .C(net12400), .Q(p2[1]) );
  DFFQX1 p2_reg_reg_0_ ( .D(N12485), .C(net12400), .Q(p2[0]) );
  DFFQX1 p2_reg_reg_2_ ( .D(N12487), .C(net12400), .Q(p2[2]) );
  DFFQX1 stop_s_reg ( .D(n1880), .C(net12400), .Q(stop) );
  DFFQX1 p2_reg_reg_6_ ( .D(N12491), .C(net12400), .Q(p2[6]) );
  DFFQX1 p2_reg_reg_3_ ( .D(N12488), .C(net12400), .Q(p2[3]) );
  DFFQX1 idle_s_reg ( .D(n1879), .C(net12400), .Q(idle) );
  DFFQX1 temp2_reg_7_ ( .D(N12730), .C(net12400), .Q(temp2_comb[7]) );
  DFFQX1 rn_reg_reg_3__7_ ( .D(n402), .C(net12521), .Q(rn_reg[231]) );
  DFFQX1 rn_reg_reg_3__2_ ( .D(n417), .C(net12521), .Q(rn_reg[226]) );
  DFFQX1 rn_reg_reg_7__7_ ( .D(n402), .C(net12541), .Q(rn_reg[199]) );
  DFFQX1 rn_reg_reg_7__2_ ( .D(n417), .C(net12541), .Q(rn_reg[194]) );
  DFFQX1 rn_reg_reg_7__6_ ( .D(n405), .C(net12541), .Q(rn_reg[198]) );
  DFFQX1 rn_reg_reg_3__6_ ( .D(n405), .C(net12521), .Q(rn_reg[230]) );
  DFFQX1 rn_reg_reg_19__7_ ( .D(n403), .C(net12601), .Q(rn_reg[103]) );
  DFFQX1 rn_reg_reg_19__6_ ( .D(n406), .C(net12601), .Q(rn_reg[102]) );
  DFFQX1 rn_reg_reg_19__2_ ( .D(n418), .C(net12601), .Q(rn_reg[98]) );
  DFFQX1 rn_reg_reg_23__7_ ( .D(n403), .C(net12621), .Q(rn_reg[71]) );
  DFFQX1 rn_reg_reg_23__6_ ( .D(n406), .C(net12621), .Q(rn_reg[70]) );
  DFFQX1 rn_reg_reg_23__2_ ( .D(n418), .C(net12621), .Q(rn_reg[66]) );
  DFFQX1 dpc_tab_reg_3__2_ ( .D(n418), .C(net12476), .Q(dpc_tab[20]) );
  DFFQX1 dpc_tab_reg_3__0_ ( .D(n426), .C(net12476), .Q(dpc_tab[18]) );
  DFFQX1 dpc_tab_reg_7__4_ ( .D(N12691), .C(net12456), .Q(dpc_tab[46]) );
  DFFQX1 dpc_tab_reg_7__2_ ( .D(n419), .C(net12456), .Q(dpc_tab[44]) );
  DFFQX1 dpc_tab_reg_7__0_ ( .D(n427), .C(net12456), .Q(dpc_tab[42]) );
  DFFQX1 rn_reg_reg_27__7_ ( .D(n403), .C(net12641), .Q(rn_reg[39]) );
  DFFQX1 rn_reg_reg_27__6_ ( .D(n407), .C(net12641), .Q(rn_reg[38]) );
  DFFQX1 rn_reg_reg_27__2_ ( .D(n419), .C(net12641), .Q(rn_reg[34]) );
  DFFQX1 rn_reg_reg_31__7_ ( .D(n404), .C(net12661), .Q(rn_reg[7]) );
  DFFQX1 rn_reg_reg_31__6_ ( .D(n407), .C(net12661), .Q(rn_reg[6]) );
  DFFQX1 rn_reg_reg_31__2_ ( .D(n420), .C(net12661), .Q(rn_reg[2]) );
  DFFQX1 rn_reg_reg_11__7_ ( .D(n404), .C(net12561), .Q(rn_reg[167]) );
  DFFQX1 rn_reg_reg_11__6_ ( .D(n407), .C(net12561), .Q(rn_reg[166]) );
  DFFQX1 rn_reg_reg_11__2_ ( .D(n420), .C(net12561), .Q(rn_reg[162]) );
  DFFQX1 rn_reg_reg_15__7_ ( .D(n1930), .C(net12581), .Q(rn_reg[135]) );
  DFFQX1 rn_reg_reg_15__6_ ( .D(n1931), .C(net12581), .Q(rn_reg[134]) );
  DFFQX1 rn_reg_reg_15__2_ ( .D(n1935), .C(net12581), .Q(rn_reg[130]) );
  DFFQX1 rn_reg_reg_0__7_ ( .D(n402), .C(net12506), .Q(rn_reg[255]) );
  DFFQX1 rn_reg_reg_0__2_ ( .D(n417), .C(net12506), .Q(rn_reg[250]) );
  DFFQX1 rn_reg_reg_4__7_ ( .D(n402), .C(net12526), .Q(rn_reg[223]) );
  DFFQX1 rn_reg_reg_4__2_ ( .D(n417), .C(net12526), .Q(rn_reg[218]) );
  DFFQX1 rn_reg_reg_0__6_ ( .D(n405), .C(net12506), .Q(rn_reg[254]) );
  DFFQX1 rn_reg_reg_4__6_ ( .D(n405), .C(net12526), .Q(rn_reg[222]) );
  DFFQX1 rn_reg_reg_16__7_ ( .D(n402), .C(net12586), .Q(rn_reg[127]) );
  DFFQX1 rn_reg_reg_16__6_ ( .D(n405), .C(net12586), .Q(rn_reg[126]) );
  DFFQX1 rn_reg_reg_16__2_ ( .D(n417), .C(net12586), .Q(rn_reg[122]) );
  DFFQX1 rn_reg_reg_20__7_ ( .D(n403), .C(net12606), .Q(rn_reg[95]) );
  DFFQX1 rn_reg_reg_20__6_ ( .D(n406), .C(net12606), .Q(rn_reg[94]) );
  DFFQX1 rn_reg_reg_20__2_ ( .D(n418), .C(net12606), .Q(rn_reg[90]) );
  DFFQX1 dpc_tab_reg_0__2_ ( .D(n419), .C(net12491), .Q(dpc_tab[2]) );
  DFFQX1 dpc_tab_reg_0__0_ ( .D(n427), .C(net12491), .Q(dpc_tab[0]) );
  DFFQX1 dpc_tab_reg_4__4_ ( .D(n413), .C(net12471), .Q(dpc_tab[28]) );
  DFFQX1 dpc_tab_reg_4__2_ ( .D(n419), .C(net12471), .Q(dpc_tab[26]) );
  DFFQX1 dpc_tab_reg_4__0_ ( .D(n427), .C(net12471), .Q(dpc_tab[24]) );
  DFFQX1 rn_reg_reg_24__7_ ( .D(n403), .C(net12626), .Q(rn_reg[63]) );
  DFFQX1 rn_reg_reg_24__6_ ( .D(n406), .C(net12626), .Q(rn_reg[62]) );
  DFFQX1 rn_reg_reg_24__2_ ( .D(n419), .C(net12626), .Q(rn_reg[58]) );
  DFFQX1 rn_reg_reg_28__7_ ( .D(n404), .C(net12646), .Q(rn_reg[31]) );
  DFFQX1 rn_reg_reg_28__6_ ( .D(n407), .C(net12646), .Q(rn_reg[30]) );
  DFFQX1 rn_reg_reg_28__2_ ( .D(n419), .C(net12646), .Q(rn_reg[26]) );
  DFFQX1 rn_reg_reg_8__7_ ( .D(n404), .C(net12546), .Q(rn_reg[191]) );
  DFFQX1 rn_reg_reg_8__6_ ( .D(n407), .C(net12546), .Q(rn_reg[190]) );
  DFFQX1 rn_reg_reg_8__2_ ( .D(n420), .C(net12546), .Q(rn_reg[186]) );
  DFFQX1 rn_reg_reg_12__7_ ( .D(n404), .C(net12566), .Q(rn_reg[159]) );
  DFFQX1 rn_reg_reg_12__6_ ( .D(n407), .C(net12566), .Q(rn_reg[158]) );
  DFFQX1 rn_reg_reg_12__2_ ( .D(n420), .C(net12566), .Q(rn_reg[154]) );
  DFFQX1 rn_reg_reg_1__7_ ( .D(n402), .C(net12511), .Q(rn_reg[247]) );
  DFFQX1 rn_reg_reg_1__2_ ( .D(n417), .C(net12511), .Q(rn_reg[242]) );
  DFFQX1 rn_reg_reg_5__7_ ( .D(n402), .C(net12531), .Q(rn_reg[215]) );
  DFFQX1 rn_reg_reg_5__2_ ( .D(n417), .C(net12531), .Q(rn_reg[210]) );
  DFFQX1 rn_reg_reg_5__6_ ( .D(n405), .C(net12531), .Q(rn_reg[214]) );
  DFFQX1 rn_reg_reg_1__6_ ( .D(n405), .C(net12511), .Q(rn_reg[246]) );
  DFFQX1 rn_reg_reg_17__7_ ( .D(n402), .C(net12591), .Q(rn_reg[119]) );
  DFFQX1 rn_reg_reg_17__6_ ( .D(n406), .C(net12591), .Q(rn_reg[118]) );
  DFFQX1 rn_reg_reg_17__2_ ( .D(n418), .C(net12591), .Q(rn_reg[114]) );
  DFFQX1 rn_reg_reg_21__7_ ( .D(n403), .C(net12611), .Q(rn_reg[87]) );
  DFFQX1 rn_reg_reg_21__6_ ( .D(n406), .C(net12611), .Q(rn_reg[86]) );
  DFFQX1 rn_reg_reg_21__2_ ( .D(n418), .C(net12611), .Q(rn_reg[82]) );
  DFFQX1 dpc_tab_reg_1__4_ ( .D(n412), .C(net12486), .Q(dpc_tab[10]) );
  DFFQX1 dpc_tab_reg_1__2_ ( .D(n418), .C(net12486), .Q(dpc_tab[8]) );
  DFFQX1 dpc_tab_reg_1__0_ ( .D(n426), .C(net12486), .Q(dpc_tab[6]) );
  DFFQX1 dpc_tab_reg_5__5_ ( .D(N12692), .C(net12466), .Q(dpc_tab[35]) );
  DFFQX1 dpc_tab_reg_5__4_ ( .D(n412), .C(net12466), .Q(dpc_tab[34]) );
  DFFQX1 dpc_tab_reg_5__2_ ( .D(n419), .C(net12466), .Q(dpc_tab[32]) );
  DFFQX1 dpc_tab_reg_5__0_ ( .D(n427), .C(net12466), .Q(dpc_tab[30]) );
  DFFQX1 rn_reg_reg_25__7_ ( .D(n403), .C(net12631), .Q(rn_reg[55]) );
  DFFQX1 rn_reg_reg_25__2_ ( .D(n419), .C(net12631), .Q(rn_reg[50]) );
  DFFQX1 rn_reg_reg_29__7_ ( .D(n404), .C(net12651), .Q(rn_reg[23]) );
  DFFQX1 rn_reg_reg_29__6_ ( .D(n407), .C(net12651), .Q(rn_reg[22]) );
  DFFQX1 rn_reg_reg_29__2_ ( .D(n420), .C(net12651), .Q(rn_reg[18]) );
  DFFQX1 rn_reg_reg_9__7_ ( .D(n404), .C(net12551), .Q(rn_reg[183]) );
  DFFQX1 rn_reg_reg_9__6_ ( .D(n407), .C(net12551), .Q(rn_reg[182]) );
  DFFQX1 rn_reg_reg_9__2_ ( .D(n420), .C(net12551), .Q(rn_reg[178]) );
  DFFQX1 rn_reg_reg_13__7_ ( .D(n404), .C(net12571), .Q(rn_reg[151]) );
  DFFQX1 rn_reg_reg_13__6_ ( .D(n1931), .C(net12571), .Q(rn_reg[150]) );
  DFFQX1 rn_reg_reg_13__2_ ( .D(n420), .C(net12571), .Q(rn_reg[146]) );
  DFFQX1 rn_reg_reg_2__7_ ( .D(n402), .C(net12516), .Q(rn_reg[239]) );
  DFFQX1 rn_reg_reg_2__2_ ( .D(n417), .C(net12516), .Q(rn_reg[234]) );
  DFFQX1 rn_reg_reg_6__7_ ( .D(n402), .C(net12536), .Q(rn_reg[207]) );
  DFFQX1 rn_reg_reg_6__2_ ( .D(n417), .C(net12536), .Q(rn_reg[202]) );
  DFFQX1 rn_reg_reg_2__6_ ( .D(n405), .C(net12516), .Q(rn_reg[238]) );
  DFFQX1 rn_reg_reg_6__6_ ( .D(n405), .C(net12536), .Q(rn_reg[206]) );
  DFFQX1 rn_reg_reg_18__7_ ( .D(n403), .C(net12596), .Q(rn_reg[111]) );
  DFFQX1 rn_reg_reg_18__6_ ( .D(n406), .C(net12596), .Q(rn_reg[110]) );
  DFFQX1 rn_reg_reg_18__2_ ( .D(n418), .C(net12596), .Q(rn_reg[106]) );
  DFFQX1 rn_reg_reg_22__7_ ( .D(n403), .C(net12616), .Q(rn_reg[79]) );
  DFFQX1 rn_reg_reg_22__6_ ( .D(n406), .C(net12616), .Q(rn_reg[78]) );
  DFFQX1 rn_reg_reg_22__2_ ( .D(n418), .C(net12616), .Q(rn_reg[74]) );
  DFFQX1 dpc_tab_reg_2__2_ ( .D(n418), .C(net12481), .Q(dpc_tab[14]) );
  DFFQX1 dpc_tab_reg_2__0_ ( .D(n426), .C(net12481), .Q(dpc_tab[12]) );
  DFFQX1 dpc_tab_reg_6__4_ ( .D(N12691), .C(net12461), .Q(dpc_tab[40]) );
  DFFQX1 dpc_tab_reg_6__2_ ( .D(n419), .C(net12461), .Q(dpc_tab[38]) );
  DFFQX1 dpc_tab_reg_6__0_ ( .D(n427), .C(net12461), .Q(dpc_tab[36]) );
  DFFQX1 rn_reg_reg_26__7_ ( .D(n403), .C(net12636), .Q(rn_reg[47]) );
  DFFQX1 rn_reg_reg_26__6_ ( .D(n406), .C(net12636), .Q(rn_reg[46]) );
  DFFQX1 rn_reg_reg_26__2_ ( .D(n419), .C(net12636), .Q(rn_reg[42]) );
  DFFQX1 rn_reg_reg_30__7_ ( .D(n404), .C(net12656), .Q(rn_reg[15]) );
  DFFQX1 rn_reg_reg_30__6_ ( .D(n407), .C(net12656), .Q(rn_reg[14]) );
  DFFQX1 rn_reg_reg_30__2_ ( .D(n420), .C(net12656), .Q(rn_reg[10]) );
  DFFQX1 rn_reg_reg_10__7_ ( .D(n404), .C(net12556), .Q(rn_reg[175]) );
  DFFQX1 rn_reg_reg_10__6_ ( .D(n407), .C(net12556), .Q(rn_reg[174]) );
  DFFQX1 rn_reg_reg_10__2_ ( .D(n420), .C(net12556), .Q(rn_reg[170]) );
  DFFQX1 rn_reg_reg_14__7_ ( .D(n1930), .C(net12576), .Q(rn_reg[143]) );
  DFFQX1 rn_reg_reg_14__6_ ( .D(n1931), .C(net12576), .Q(rn_reg[142]) );
  DFFQX1 rn_reg_reg_14__2_ ( .D(n420), .C(net12576), .Q(rn_reg[138]) );
  DFFQX1 dec_cop_reg_7_ ( .D(N10589), .C(net12400), .Q(dec_cop[7]) );
  DFFQX1 sp_reg_reg_5_ ( .D(N12702), .C(net12400), .Q(sp[5]) );
  DFFQX1 f1_reg ( .D(n1883), .C(net12400), .Q(f1) );
  DFFQX1 sp_reg_reg_6_ ( .D(N12703), .C(net12400), .Q(sp[6]) );
  DFFQX1 dph_reg_reg_3__6_ ( .D(N12527), .C(net12436), .Q(dph_reg[30]) );
  DFFQX1 dph_reg_reg_3__5_ ( .D(N12526), .C(net12436), .Q(dph_reg[29]) );
  DFFQX1 dph_reg_reg_3__4_ ( .D(N12525), .C(net12436), .Q(dph_reg[28]) );
  DFFQX1 dph_reg_reg_3__3_ ( .D(N12524), .C(net12436), .Q(dph_reg[27]) );
  DFFQX1 dph_reg_reg_3__2_ ( .D(N12523), .C(net12436), .Q(dph_reg[26]) );
  DFFQX1 dph_reg_reg_3__1_ ( .D(N12522), .C(net12436), .Q(dph_reg[25]) );
  DFFQX1 dpl_reg_reg_3__5_ ( .D(N12598), .C(net12436), .Q(dpl_reg[29]) );
  DFFQX1 dpl_reg_reg_3__4_ ( .D(N12597), .C(net12436), .Q(dpl_reg[28]) );
  DFFQX1 dpl_reg_reg_3__2_ ( .D(N12595), .C(net12436), .Q(dpl_reg[26]) );
  DFFQX1 dph_reg_reg_7__6_ ( .D(N12563), .C(net12416), .Q(dph_reg[62]) );
  DFFQX1 dph_reg_reg_7__5_ ( .D(N12562), .C(net12416), .Q(dph_reg[61]) );
  DFFQX1 dph_reg_reg_7__4_ ( .D(N12561), .C(net12416), .Q(dph_reg[60]) );
  DFFQX1 dph_reg_reg_7__2_ ( .D(N12559), .C(net12416), .Q(dph_reg[58]) );
  DFFQX1 dpl_reg_reg_7__5_ ( .D(N12634), .C(net12416), .Q(dpl_reg[61]) );
  DFFQX1 dpl_reg_reg_7__4_ ( .D(N12633), .C(net12416), .Q(dpl_reg[60]) );
  DFFQX1 dpl_reg_reg_7__3_ ( .D(N12632), .C(net12416), .Q(dpl_reg[59]) );
  DFFQX1 dpl_reg_reg_7__2_ ( .D(N12631), .C(net12416), .Q(dpl_reg[58]) );
  DFFQX1 dph_reg_reg_7__0_ ( .D(N12557), .C(net12416), .Q(dph_reg[56]) );
  DFFQX1 dph_reg_reg_3__0_ ( .D(N12521), .C(net12436), .Q(dph_reg[24]) );
  DFFQX1 dph_reg_reg_0__6_ ( .D(N12500), .C(net12451), .Q(dph_reg[6]) );
  DFFQX1 dph_reg_reg_0__5_ ( .D(N12499), .C(net12451), .Q(dph_reg[5]) );
  DFFQX1 dph_reg_reg_0__4_ ( .D(N12498), .C(net12451), .Q(dph_reg[4]) );
  DFFQX1 dph_reg_reg_0__2_ ( .D(N12496), .C(net12451), .Q(dph_reg[2]) );
  DFFQX1 dpl_reg_reg_0__5_ ( .D(N12571), .C(net12451), .Q(dpl_reg[5]) );
  DFFQX1 dpl_reg_reg_0__4_ ( .D(N12570), .C(net12451), .Q(dpl_reg[4]) );
  DFFQX1 dpl_reg_reg_0__2_ ( .D(N12568), .C(net12451), .Q(dpl_reg[2]) );
  DFFQX1 dph_reg_reg_4__6_ ( .D(N12536), .C(net12431), .Q(dph_reg[38]) );
  DFFQX1 dph_reg_reg_4__5_ ( .D(N12535), .C(net12431), .Q(dph_reg[37]) );
  DFFQX1 dph_reg_reg_4__4_ ( .D(N12534), .C(net12431), .Q(dph_reg[36]) );
  DFFQX1 dph_reg_reg_4__2_ ( .D(N12532), .C(net12431), .Q(dph_reg[34]) );
  DFFQX1 dpl_reg_reg_4__5_ ( .D(N12607), .C(net12431), .Q(dpl_reg[37]) );
  DFFQX1 dpl_reg_reg_4__4_ ( .D(N12606), .C(net12431), .Q(dpl_reg[36]) );
  DFFQX1 dpl_reg_reg_4__3_ ( .D(N12605), .C(net12431), .Q(dpl_reg[35]) );
  DFFQX1 dpl_reg_reg_4__2_ ( .D(N12604), .C(net12431), .Q(dpl_reg[34]) );
  DFFQX1 dph_reg_reg_4__0_ ( .D(N12530), .C(net12431), .Q(dph_reg[32]) );
  DFFQX1 dph_reg_reg_0__0_ ( .D(N12494), .C(net12451), .Q(dph_reg[0]) );
  DFFQX1 dph_reg_reg_1__6_ ( .D(N12509), .C(net12446), .Q(dph_reg[14]) );
  DFFQX1 dph_reg_reg_1__5_ ( .D(N12508), .C(net12446), .Q(dph_reg[13]) );
  DFFQX1 dph_reg_reg_1__4_ ( .D(N12507), .C(net12446), .Q(dph_reg[12]) );
  DFFQX1 dph_reg_reg_1__2_ ( .D(N12505), .C(net12446), .Q(dph_reg[10]) );
  DFFQX1 dpl_reg_reg_1__5_ ( .D(N12580), .C(net12446), .Q(dpl_reg[13]) );
  DFFQX1 dpl_reg_reg_1__4_ ( .D(N12579), .C(net12446), .Q(dpl_reg[12]) );
  DFFQX1 dpl_reg_reg_1__3_ ( .D(N12578), .C(net12446), .Q(dpl_reg[11]) );
  DFFQX1 dpl_reg_reg_1__2_ ( .D(N12577), .C(net12446), .Q(dpl_reg[10]) );
  DFFQX1 dph_reg_reg_5__6_ ( .D(N12545), .C(net12426), .Q(dph_reg[46]) );
  DFFQX1 dph_reg_reg_5__5_ ( .D(N12544), .C(net12426), .Q(dph_reg[45]) );
  DFFQX1 dph_reg_reg_5__4_ ( .D(N12543), .C(net12426), .Q(dph_reg[44]) );
  DFFQX1 dph_reg_reg_5__2_ ( .D(N12541), .C(net12426), .Q(dph_reg[42]) );
  DFFQX1 dpl_reg_reg_5__5_ ( .D(N12616), .C(net12426), .Q(dpl_reg[45]) );
  DFFQX1 dpl_reg_reg_5__4_ ( .D(N12615), .C(net12426), .Q(dpl_reg[44]) );
  DFFQX1 dpl_reg_reg_5__3_ ( .D(N12614), .C(net12426), .Q(dpl_reg[43]) );
  DFFQX1 dpl_reg_reg_5__2_ ( .D(N12613), .C(net12426), .Q(dpl_reg[42]) );
  DFFQX1 dph_reg_reg_5__0_ ( .D(N12539), .C(net12426), .Q(dph_reg[40]) );
  DFFQX1 dph_reg_reg_1__0_ ( .D(N12503), .C(net12446), .Q(dph_reg[8]) );
  DFFQX1 dph_reg_reg_2__6_ ( .D(N12518), .C(net12441), .Q(dph_reg[22]) );
  DFFQX1 dph_reg_reg_2__5_ ( .D(N12517), .C(net12441), .Q(dph_reg[21]) );
  DFFQX1 dph_reg_reg_2__4_ ( .D(N12516), .C(net12441), .Q(dph_reg[20]) );
  DFFQX1 dph_reg_reg_2__3_ ( .D(N12515), .C(net12441), .Q(dph_reg[19]) );
  DFFQX1 dph_reg_reg_2__2_ ( .D(N12514), .C(net12441), .Q(dph_reg[18]) );
  DFFQX1 dph_reg_reg_2__1_ ( .D(N12513), .C(net12441), .Q(dph_reg[17]) );
  DFFQX1 dpl_reg_reg_2__5_ ( .D(N12589), .C(net12441), .Q(dpl_reg[21]) );
  DFFQX1 dpl_reg_reg_2__4_ ( .D(N12588), .C(net12441), .Q(dpl_reg[20]) );
  DFFQX1 dpl_reg_reg_2__2_ ( .D(N12586), .C(net12441), .Q(dpl_reg[18]) );
  DFFQX1 dph_reg_reg_6__6_ ( .D(N12554), .C(net12421), .Q(dph_reg[54]) );
  DFFQX1 dph_reg_reg_6__5_ ( .D(N12553), .C(net12421), .Q(dph_reg[53]) );
  DFFQX1 dph_reg_reg_6__4_ ( .D(N12552), .C(net12421), .Q(dph_reg[52]) );
  DFFQX1 dph_reg_reg_6__2_ ( .D(N12550), .C(net12421), .Q(dph_reg[50]) );
  DFFQX1 dpl_reg_reg_6__5_ ( .D(N12625), .C(net12421), .Q(dpl_reg[53]) );
  DFFQX1 dpl_reg_reg_6__4_ ( .D(N12624), .C(net12421), .Q(dpl_reg[52]) );
  DFFQX1 dpl_reg_reg_6__3_ ( .D(N12623), .C(net12421), .Q(dpl_reg[51]) );
  DFFQX1 dpl_reg_reg_6__2_ ( .D(N12622), .C(net12421), .Q(dpl_reg[50]) );
  DFFQX1 dph_reg_reg_6__0_ ( .D(N12548), .C(net12421), .Q(dph_reg[48]) );
  DFFQX1 dph_reg_reg_2__0_ ( .D(N12512), .C(net12441), .Q(dph_reg[16]) );
  DFFQX1 dec_cop_reg_6_ ( .D(N10588), .C(net12400), .Q(dec_cop[6]) );
  DFFQX1 multempreg_reg_0_ ( .D(N13325), .C(net12666), .Q(multempreg[0]) );
  DFFQX1 ckcon_r_reg_7_ ( .D(N12972), .C(net12400), .Q(ckcon[7]) );
  DFFQX1 rmwinstr_reg ( .D(N690), .C(net12400), .Q(rmwinstr) );
  DFFQX1 bitno_reg_2_ ( .D(N11494), .C(net12411), .Q(N345) );
  DFFQX1 ramdatao_r_reg_6_ ( .D(N11504), .C(net12400), .Q(ramdatao[6]) );
  DFFQX1 ramdatao_r_reg_5_ ( .D(N11503), .C(net12400), .Q(ramdatao[5]) );
  DFFQX1 ramdatao_r_reg_7_ ( .D(N11505), .C(net12400), .Q(ramdatao[7]) );
  DFFQX1 rn_reg_reg_3__3_ ( .D(n414), .C(net12521), .Q(rn_reg[227]) );
  DFFQX1 rn_reg_reg_3__1_ ( .D(n421), .C(net12521), .Q(rn_reg[225]) );
  DFFQX1 rn_reg_reg_3__0_ ( .D(n425), .C(net12521), .Q(rn_reg[224]) );
  DFFQX1 rn_reg_reg_7__3_ ( .D(n414), .C(net12541), .Q(rn_reg[195]) );
  DFFQX1 rn_reg_reg_7__1_ ( .D(n421), .C(net12541), .Q(rn_reg[193]) );
  DFFQX1 rn_reg_reg_7__0_ ( .D(n425), .C(net12541), .Q(rn_reg[192]) );
  DFFQX1 rn_reg_reg_7__4_ ( .D(n411), .C(net12541), .Q(rn_reg[196]) );
  DFFQX1 rn_reg_reg_3__4_ ( .D(n411), .C(net12521), .Q(rn_reg[228]) );
  DFFQX1 rn_reg_reg_7__5_ ( .D(n408), .C(net12541), .Q(rn_reg[197]) );
  DFFQX1 rn_reg_reg_3__5_ ( .D(n408), .C(net12521), .Q(rn_reg[229]) );
  DFFQX1 rn_reg_reg_19__5_ ( .D(n409), .C(net12601), .Q(rn_reg[101]) );
  DFFQX1 rn_reg_reg_19__4_ ( .D(n412), .C(net12601), .Q(rn_reg[100]) );
  DFFQX1 rn_reg_reg_19__1_ ( .D(n422), .C(net12601), .Q(rn_reg[97]) );
  DFFQX1 rn_reg_reg_19__0_ ( .D(n426), .C(net12601), .Q(rn_reg[96]) );
  DFFQX1 rn_reg_reg_23__5_ ( .D(n409), .C(net12621), .Q(rn_reg[69]) );
  DFFQX1 rn_reg_reg_23__4_ ( .D(n412), .C(net12621), .Q(rn_reg[68]) );
  DFFQX1 rn_reg_reg_23__3_ ( .D(n415), .C(net12621), .Q(rn_reg[67]) );
  DFFQX1 rn_reg_reg_23__1_ ( .D(n422), .C(net12621), .Q(rn_reg[65]) );
  DFFQX1 rn_reg_reg_23__0_ ( .D(n426), .C(net12621), .Q(rn_reg[64]) );
  DFFQX1 dpc_tab_reg_3__3_ ( .D(N12690), .C(net12476), .Q(dpc_tab[21]) );
  DFFQX1 dpc_tab_reg_3__1_ ( .D(n422), .C(net12476), .Q(dpc_tab[19]) );
  DFFQX1 dpc_tab_reg_7__3_ ( .D(N12690), .C(net12456), .Q(dpc_tab[45]) );
  DFFQX1 dpc_tab_reg_7__1_ ( .D(n423), .C(net12456), .Q(dpc_tab[43]) );
  DFFQX1 rn_reg_reg_27__5_ ( .D(n410), .C(net12641), .Q(rn_reg[37]) );
  DFFQX1 rn_reg_reg_27__4_ ( .D(n413), .C(net12641), .Q(rn_reg[36]) );
  DFFQX1 rn_reg_reg_27__1_ ( .D(n423), .C(net12641), .Q(rn_reg[33]) );
  DFFQX1 rn_reg_reg_27__0_ ( .D(n427), .C(net12641), .Q(rn_reg[32]) );
  DFFQX1 rn_reg_reg_31__5_ ( .D(n410), .C(net12661), .Q(rn_reg[5]) );
  DFFQX1 rn_reg_reg_31__4_ ( .D(n413), .C(net12661), .Q(rn_reg[4]) );
  DFFQX1 rn_reg_reg_31__3_ ( .D(n416), .C(net12661), .Q(rn_reg[3]) );
  DFFQX1 rn_reg_reg_31__1_ ( .D(n424), .C(net12661), .Q(rn_reg[1]) );
  DFFQX1 rn_reg_reg_31__0_ ( .D(n428), .C(net12661), .Q(rn_reg[0]) );
  DFFQX1 rn_reg_reg_11__5_ ( .D(n1932), .C(net12561), .Q(rn_reg[165]) );
  DFFQX1 rn_reg_reg_11__4_ ( .D(n1933), .C(net12561), .Q(rn_reg[164]) );
  DFFQX1 rn_reg_reg_11__3_ ( .D(n1934), .C(net12561), .Q(rn_reg[163]) );
  DFFQX1 rn_reg_reg_11__1_ ( .D(n424), .C(net12561), .Q(rn_reg[161]) );
  DFFQX1 rn_reg_reg_11__0_ ( .D(n428), .C(net12561), .Q(rn_reg[160]) );
  DFFQX1 rn_reg_reg_15__5_ ( .D(n1932), .C(net12581), .Q(rn_reg[133]) );
  DFFQX1 rn_reg_reg_15__4_ ( .D(n1933), .C(net12581), .Q(rn_reg[132]) );
  DFFQX1 rn_reg_reg_15__3_ ( .D(n1934), .C(net12581), .Q(rn_reg[131]) );
  DFFQX1 rn_reg_reg_15__1_ ( .D(n1936), .C(net12581), .Q(rn_reg[129]) );
  DFFQX1 rn_reg_reg_15__0_ ( .D(n1937), .C(net12581), .Q(rn_reg[128]) );
  DFFQX1 rn_reg_reg_0__3_ ( .D(n414), .C(net12506), .Q(rn_reg[251]) );
  DFFQX1 rn_reg_reg_0__1_ ( .D(n421), .C(net12506), .Q(rn_reg[249]) );
  DFFQX1 rn_reg_reg_0__0_ ( .D(n425), .C(net12506), .Q(rn_reg[248]) );
  DFFQX1 rn_reg_reg_4__3_ ( .D(n414), .C(net12526), .Q(rn_reg[219]) );
  DFFQX1 rn_reg_reg_4__1_ ( .D(n421), .C(net12526), .Q(rn_reg[217]) );
  DFFQX1 rn_reg_reg_4__0_ ( .D(n425), .C(net12526), .Q(rn_reg[216]) );
  DFFQX1 rn_reg_reg_0__4_ ( .D(n411), .C(net12506), .Q(rn_reg[252]) );
  DFFQX1 rn_reg_reg_4__4_ ( .D(n411), .C(net12526), .Q(rn_reg[220]) );
  DFFQX1 rn_reg_reg_0__5_ ( .D(n408), .C(net12506), .Q(rn_reg[253]) );
  DFFQX1 rn_reg_reg_4__5_ ( .D(n408), .C(net12526), .Q(rn_reg[221]) );
  DFFQX1 rn_reg_reg_16__5_ ( .D(n408), .C(net12586), .Q(rn_reg[125]) );
  DFFQX1 rn_reg_reg_16__4_ ( .D(n411), .C(net12586), .Q(rn_reg[124]) );
  DFFQX1 rn_reg_reg_16__1_ ( .D(n421), .C(net12586), .Q(rn_reg[121]) );
  DFFQX1 rn_reg_reg_16__0_ ( .D(n425), .C(net12586), .Q(rn_reg[120]) );
  DFFQX1 rn_reg_reg_20__5_ ( .D(n409), .C(net12606), .Q(rn_reg[93]) );
  DFFQX1 rn_reg_reg_20__4_ ( .D(n412), .C(net12606), .Q(rn_reg[92]) );
  DFFQX1 rn_reg_reg_20__1_ ( .D(n422), .C(net12606), .Q(rn_reg[89]) );
  DFFQX1 rn_reg_reg_20__0_ ( .D(n426), .C(net12606), .Q(rn_reg[88]) );
  DFFQX1 dpc_tab_reg_0__3_ ( .D(n415), .C(net12491), .Q(dpc_tab[3]) );
  DFFQX1 dpc_tab_reg_0__1_ ( .D(n423), .C(net12491), .Q(dpc_tab[1]) );
  DFFQX1 dpc_tab_reg_4__3_ ( .D(n416), .C(net12471), .Q(dpc_tab[27]) );
  DFFQX1 dpc_tab_reg_4__1_ ( .D(n423), .C(net12471), .Q(dpc_tab[25]) );
  DFFQX1 rn_reg_reg_24__5_ ( .D(n410), .C(net12626), .Q(rn_reg[61]) );
  DFFQX1 rn_reg_reg_24__4_ ( .D(n413), .C(net12626), .Q(rn_reg[60]) );
  DFFQX1 rn_reg_reg_24__1_ ( .D(n423), .C(net12626), .Q(rn_reg[57]) );
  DFFQX1 rn_reg_reg_24__0_ ( .D(n427), .C(net12626), .Q(rn_reg[56]) );
  DFFQX1 rn_reg_reg_28__5_ ( .D(n410), .C(net12646), .Q(rn_reg[29]) );
  DFFQX1 rn_reg_reg_28__4_ ( .D(n413), .C(net12646), .Q(rn_reg[28]) );
  DFFQX1 rn_reg_reg_28__1_ ( .D(n423), .C(net12646), .Q(rn_reg[25]) );
  DFFQX1 rn_reg_reg_28__0_ ( .D(n427), .C(net12646), .Q(rn_reg[24]) );
  DFFQX1 rn_reg_reg_8__5_ ( .D(n410), .C(net12546), .Q(rn_reg[189]) );
  DFFQX1 rn_reg_reg_8__4_ ( .D(n413), .C(net12546), .Q(rn_reg[188]) );
  DFFQX1 rn_reg_reg_8__3_ ( .D(n416), .C(net12546), .Q(rn_reg[187]) );
  DFFQX1 rn_reg_reg_8__1_ ( .D(n424), .C(net12546), .Q(rn_reg[185]) );
  DFFQX1 rn_reg_reg_8__0_ ( .D(n428), .C(net12546), .Q(rn_reg[184]) );
  DFFQX1 rn_reg_reg_12__5_ ( .D(n1932), .C(net12566), .Q(rn_reg[157]) );
  DFFQX1 rn_reg_reg_12__4_ ( .D(n1933), .C(net12566), .Q(rn_reg[156]) );
  DFFQX1 rn_reg_reg_12__3_ ( .D(n1934), .C(net12566), .Q(rn_reg[155]) );
  DFFQX1 rn_reg_reg_12__1_ ( .D(n424), .C(net12566), .Q(rn_reg[153]) );
  DFFQX1 rn_reg_reg_12__0_ ( .D(n428), .C(net12566), .Q(rn_reg[152]) );
  DFFQX1 rn_reg_reg_1__3_ ( .D(n414), .C(net12511), .Q(rn_reg[243]) );
  DFFQX1 rn_reg_reg_1__1_ ( .D(n421), .C(net12511), .Q(rn_reg[241]) );
  DFFQX1 rn_reg_reg_1__0_ ( .D(n425), .C(net12511), .Q(rn_reg[240]) );
  DFFQX1 rn_reg_reg_5__3_ ( .D(n414), .C(net12531), .Q(rn_reg[211]) );
  DFFQX1 rn_reg_reg_5__1_ ( .D(n421), .C(net12531), .Q(rn_reg[209]) );
  DFFQX1 rn_reg_reg_5__0_ ( .D(n425), .C(net12531), .Q(rn_reg[208]) );
  DFFQX1 rn_reg_reg_5__4_ ( .D(n411), .C(net12531), .Q(rn_reg[212]) );
  DFFQX1 rn_reg_reg_1__4_ ( .D(n411), .C(net12511), .Q(rn_reg[244]) );
  DFFQX1 rn_reg_reg_5__5_ ( .D(n408), .C(net12531), .Q(rn_reg[213]) );
  DFFQX1 rn_reg_reg_1__5_ ( .D(n408), .C(net12511), .Q(rn_reg[245]) );
  DFFQX1 rn_reg_reg_17__5_ ( .D(n409), .C(net12591), .Q(rn_reg[117]) );
  DFFQX1 rn_reg_reg_17__4_ ( .D(n412), .C(net12591), .Q(rn_reg[116]) );
  DFFQX1 rn_reg_reg_17__1_ ( .D(n422), .C(net12591), .Q(rn_reg[113]) );
  DFFQX1 rn_reg_reg_17__0_ ( .D(n426), .C(net12591), .Q(rn_reg[112]) );
  DFFQX1 rn_reg_reg_21__5_ ( .D(n409), .C(net12611), .Q(rn_reg[85]) );
  DFFQX1 rn_reg_reg_21__4_ ( .D(n412), .C(net12611), .Q(rn_reg[84]) );
  DFFQX1 rn_reg_reg_21__1_ ( .D(n422), .C(net12611), .Q(rn_reg[81]) );
  DFFQX1 rn_reg_reg_21__0_ ( .D(n426), .C(net12611), .Q(rn_reg[80]) );
  DFFQX1 dpc_tab_reg_1__3_ ( .D(N12690), .C(net12486), .Q(dpc_tab[9]) );
  DFFQX1 dpc_tab_reg_1__1_ ( .D(n422), .C(net12486), .Q(dpc_tab[7]) );
  DFFQX1 dpc_tab_reg_5__3_ ( .D(N12690), .C(net12466), .Q(dpc_tab[33]) );
  DFFQX1 dpc_tab_reg_5__1_ ( .D(n423), .C(net12466), .Q(dpc_tab[31]) );
  DFFQX1 rn_reg_reg_25__6_ ( .D(n406), .C(net12631), .Q(rn_reg[54]) );
  DFFQX1 rn_reg_reg_25__5_ ( .D(n410), .C(net12631), .Q(rn_reg[53]) );
  DFFQX1 rn_reg_reg_25__4_ ( .D(n413), .C(net12631), .Q(rn_reg[52]) );
  DFFQX1 rn_reg_reg_25__1_ ( .D(n423), .C(net12631), .Q(rn_reg[49]) );
  DFFQX1 rn_reg_reg_25__0_ ( .D(n427), .C(net12631), .Q(rn_reg[48]) );
  DFFQX1 rn_reg_reg_29__5_ ( .D(n410), .C(net12651), .Q(rn_reg[21]) );
  DFFQX1 rn_reg_reg_29__4_ ( .D(n413), .C(net12651), .Q(rn_reg[20]) );
  DFFQX1 rn_reg_reg_29__1_ ( .D(n424), .C(net12651), .Q(rn_reg[17]) );
  DFFQX1 rn_reg_reg_29__0_ ( .D(n428), .C(net12651), .Q(rn_reg[16]) );
  DFFQX1 rn_reg_reg_9__5_ ( .D(n1932), .C(net12551), .Q(rn_reg[181]) );
  DFFQX1 rn_reg_reg_9__4_ ( .D(n1933), .C(net12551), .Q(rn_reg[180]) );
  DFFQX1 rn_reg_reg_9__3_ ( .D(n1934), .C(net12551), .Q(rn_reg[179]) );
  DFFQX1 rn_reg_reg_9__1_ ( .D(n424), .C(net12551), .Q(rn_reg[177]) );
  DFFQX1 rn_reg_reg_9__0_ ( .D(n428), .C(net12551), .Q(rn_reg[176]) );
  DFFQX1 rn_reg_reg_13__5_ ( .D(n1932), .C(net12571), .Q(rn_reg[149]) );
  DFFQX1 rn_reg_reg_13__4_ ( .D(n1933), .C(net12571), .Q(rn_reg[148]) );
  DFFQX1 rn_reg_reg_13__3_ ( .D(n1934), .C(net12571), .Q(rn_reg[147]) );
  DFFQX1 rn_reg_reg_13__1_ ( .D(n424), .C(net12571), .Q(rn_reg[145]) );
  DFFQX1 rn_reg_reg_13__0_ ( .D(n428), .C(net12571), .Q(rn_reg[144]) );
  DFFQX1 rn_reg_reg_2__3_ ( .D(n414), .C(net12516), .Q(rn_reg[235]) );
  DFFQX1 rn_reg_reg_2__1_ ( .D(n421), .C(net12516), .Q(rn_reg[233]) );
  DFFQX1 rn_reg_reg_2__0_ ( .D(n425), .C(net12516), .Q(rn_reg[232]) );
  DFFQX1 rn_reg_reg_6__3_ ( .D(n414), .C(net12536), .Q(rn_reg[203]) );
  DFFQX1 rn_reg_reg_6__1_ ( .D(n421), .C(net12536), .Q(rn_reg[201]) );
  DFFQX1 rn_reg_reg_6__0_ ( .D(n425), .C(net12536), .Q(rn_reg[200]) );
  DFFQX1 rn_reg_reg_2__4_ ( .D(n411), .C(net12516), .Q(rn_reg[236]) );
  DFFQX1 rn_reg_reg_6__4_ ( .D(n411), .C(net12536), .Q(rn_reg[204]) );
  DFFQX1 rn_reg_reg_2__5_ ( .D(n408), .C(net12516), .Q(rn_reg[237]) );
  DFFQX1 rn_reg_reg_6__5_ ( .D(n408), .C(net12536), .Q(rn_reg[205]) );
  DFFQX1 rn_reg_reg_18__5_ ( .D(n409), .C(net12596), .Q(rn_reg[109]) );
  DFFQX1 rn_reg_reg_18__4_ ( .D(n412), .C(net12596), .Q(rn_reg[108]) );
  DFFQX1 rn_reg_reg_18__1_ ( .D(n422), .C(net12596), .Q(rn_reg[105]) );
  DFFQX1 rn_reg_reg_18__0_ ( .D(n426), .C(net12596), .Q(rn_reg[104]) );
  DFFQX1 rn_reg_reg_22__5_ ( .D(n409), .C(net12616), .Q(rn_reg[77]) );
  DFFQX1 rn_reg_reg_22__4_ ( .D(n412), .C(net12616), .Q(rn_reg[76]) );
  DFFQX1 rn_reg_reg_22__3_ ( .D(n415), .C(net12616), .Q(rn_reg[75]) );
  DFFQX1 rn_reg_reg_22__1_ ( .D(n422), .C(net12616), .Q(rn_reg[73]) );
  DFFQX1 rn_reg_reg_22__0_ ( .D(n426), .C(net12616), .Q(rn_reg[72]) );
  DFFQX1 dpc_tab_reg_2__3_ ( .D(n415), .C(net12481), .Q(dpc_tab[15]) );
  DFFQX1 dpc_tab_reg_2__1_ ( .D(n422), .C(net12481), .Q(dpc_tab[13]) );
  DFFQX1 dpc_tab_reg_6__3_ ( .D(n415), .C(net12461), .Q(dpc_tab[39]) );
  DFFQX1 dpc_tab_reg_6__1_ ( .D(n423), .C(net12461), .Q(dpc_tab[37]) );
  DFFQX1 rn_reg_reg_26__5_ ( .D(n410), .C(net12636), .Q(rn_reg[45]) );
  DFFQX1 rn_reg_reg_26__4_ ( .D(n413), .C(net12636), .Q(rn_reg[44]) );
  DFFQX1 rn_reg_reg_26__1_ ( .D(n423), .C(net12636), .Q(rn_reg[41]) );
  DFFQX1 rn_reg_reg_26__0_ ( .D(n427), .C(net12636), .Q(rn_reg[40]) );
  DFFQX1 rn_reg_reg_30__5_ ( .D(n410), .C(net12656), .Q(rn_reg[13]) );
  DFFQX1 rn_reg_reg_30__4_ ( .D(n413), .C(net12656), .Q(rn_reg[12]) );
  DFFQX1 rn_reg_reg_30__3_ ( .D(n416), .C(net12656), .Q(rn_reg[11]) );
  DFFQX1 rn_reg_reg_30__1_ ( .D(n424), .C(net12656), .Q(rn_reg[9]) );
  DFFQX1 rn_reg_reg_30__0_ ( .D(n428), .C(net12656), .Q(rn_reg[8]) );
  DFFQX1 rn_reg_reg_10__5_ ( .D(n1932), .C(net12556), .Q(rn_reg[173]) );
  DFFQX1 rn_reg_reg_10__4_ ( .D(n1933), .C(net12556), .Q(rn_reg[172]) );
  DFFQX1 rn_reg_reg_10__3_ ( .D(n1934), .C(net12556), .Q(rn_reg[171]) );
  DFFQX1 rn_reg_reg_10__1_ ( .D(n424), .C(net12556), .Q(rn_reg[169]) );
  DFFQX1 rn_reg_reg_10__0_ ( .D(n428), .C(net12556), .Q(rn_reg[168]) );
  DFFQX1 rn_reg_reg_14__5_ ( .D(n1932), .C(net12576), .Q(rn_reg[141]) );
  DFFQX1 rn_reg_reg_14__4_ ( .D(n1933), .C(net12576), .Q(rn_reg[140]) );
  DFFQX1 rn_reg_reg_14__3_ ( .D(n1934), .C(net12576), .Q(rn_reg[139]) );
  DFFQX1 rn_reg_reg_14__1_ ( .D(n424), .C(net12576), .Q(rn_reg[137]) );
  DFFQX1 rn_reg_reg_14__0_ ( .D(n428), .C(net12576), .Q(rn_reg[136]) );
  DFFQX1 sp_reg_reg_4_ ( .D(N12701), .C(net12400), .Q(sp[4]) );
  DFFQX1 sp_reg_reg_3_ ( .D(N12700), .C(net12400), .Q(sp[3]) );
  DFFQX1 dph_reg_reg_3__7_ ( .D(N12528), .C(net12436), .Q(dph_reg[31]) );
  DFFQX1 dpl_reg_reg_3__7_ ( .D(N12600), .C(net12436), .Q(dpl_reg[31]) );
  DFFQX1 dpl_reg_reg_3__6_ ( .D(N12599), .C(net12436), .Q(dpl_reg[30]) );
  DFFQX1 dpl_reg_reg_3__1_ ( .D(N12594), .C(net12436), .Q(dpl_reg[25]) );
  DFFQX1 dpl_reg_reg_3__0_ ( .D(N12593), .C(net12436), .Q(dpl_reg[24]) );
  DFFQX1 dph_reg_reg_7__7_ ( .D(N12564), .C(net12416), .Q(dph_reg[63]) );
  DFFQX1 dph_reg_reg_7__3_ ( .D(N12560), .C(net12416), .Q(dph_reg[59]) );
  DFFQX1 dph_reg_reg_7__1_ ( .D(N12558), .C(net12416), .Q(dph_reg[57]) );
  DFFQX1 dpl_reg_reg_7__7_ ( .D(N12636), .C(net12416), .Q(dpl_reg[63]) );
  DFFQX1 dpl_reg_reg_7__6_ ( .D(N12635), .C(net12416), .Q(dpl_reg[62]) );
  DFFQX1 dpl_reg_reg_7__1_ ( .D(N12630), .C(net12416), .Q(dpl_reg[57]) );
  DFFQX1 dpl_reg_reg_7__0_ ( .D(N12629), .C(net12416), .Q(dpl_reg[56]) );
  DFFQX1 dph_reg_reg_0__7_ ( .D(N12501), .C(net12451), .Q(dph_reg[7]) );
  DFFQX1 dph_reg_reg_0__3_ ( .D(N12497), .C(net12451), .Q(dph_reg[3]) );
  DFFQX1 dph_reg_reg_0__1_ ( .D(N12495), .C(net12451), .Q(dph_reg[1]) );
  DFFQX1 dpl_reg_reg_0__7_ ( .D(N12573), .C(net12451), .Q(dpl_reg[7]) );
  DFFQX1 dpl_reg_reg_0__6_ ( .D(N12572), .C(net12451), .Q(dpl_reg[6]) );
  DFFQX1 dpl_reg_reg_0__1_ ( .D(N12567), .C(net12451), .Q(dpl_reg[1]) );
  DFFQX1 dpl_reg_reg_0__0_ ( .D(N12566), .C(net12451), .Q(dpl_reg[0]) );
  DFFQX1 dph_reg_reg_4__7_ ( .D(N12537), .C(net12431), .Q(dph_reg[39]) );
  DFFQX1 dph_reg_reg_4__3_ ( .D(N12533), .C(net12431), .Q(dph_reg[35]) );
  DFFQX1 dph_reg_reg_4__1_ ( .D(N12531), .C(net12431), .Q(dph_reg[33]) );
  DFFQX1 dpl_reg_reg_4__7_ ( .D(N12609), .C(net12431), .Q(dpl_reg[39]) );
  DFFQX1 dpl_reg_reg_4__6_ ( .D(N12608), .C(net12431), .Q(dpl_reg[38]) );
  DFFQX1 dpl_reg_reg_4__1_ ( .D(N12603), .C(net12431), .Q(dpl_reg[33]) );
  DFFQX1 dpl_reg_reg_4__0_ ( .D(N12602), .C(net12431), .Q(dpl_reg[32]) );
  DFFQX1 dph_reg_reg_1__7_ ( .D(N12510), .C(net12446), .Q(dph_reg[15]) );
  DFFQX1 dph_reg_reg_1__3_ ( .D(N12506), .C(net12446), .Q(dph_reg[11]) );
  DFFQX1 dph_reg_reg_1__1_ ( .D(N12504), .C(net12446), .Q(dph_reg[9]) );
  DFFQX1 dpl_reg_reg_1__7_ ( .D(N12582), .C(net12446), .Q(dpl_reg[15]) );
  DFFQX1 dpl_reg_reg_1__6_ ( .D(N12581), .C(net12446), .Q(dpl_reg[14]) );
  DFFQX1 dpl_reg_reg_1__1_ ( .D(N12576), .C(net12446), .Q(dpl_reg[9]) );
  DFFQX1 dpl_reg_reg_1__0_ ( .D(N12575), .C(net12446), .Q(dpl_reg[8]) );
  DFFQX1 dph_reg_reg_5__7_ ( .D(N12546), .C(net12426), .Q(dph_reg[47]) );
  DFFQX1 dph_reg_reg_5__3_ ( .D(N12542), .C(net12426), .Q(dph_reg[43]) );
  DFFQX1 dph_reg_reg_5__1_ ( .D(N12540), .C(net12426), .Q(dph_reg[41]) );
  DFFQX1 dpl_reg_reg_5__7_ ( .D(N12618), .C(net12426), .Q(dpl_reg[47]) );
  DFFQX1 dpl_reg_reg_5__6_ ( .D(N12617), .C(net12426), .Q(dpl_reg[46]) );
  DFFQX1 dpl_reg_reg_5__1_ ( .D(N12612), .C(net12426), .Q(dpl_reg[41]) );
  DFFQX1 dpl_reg_reg_5__0_ ( .D(N12611), .C(net12426), .Q(dpl_reg[40]) );
  DFFQX1 dph_reg_reg_2__7_ ( .D(N12519), .C(net12441), .Q(dph_reg[23]) );
  DFFQX1 dpl_reg_reg_2__7_ ( .D(N12591), .C(net12441), .Q(dpl_reg[23]) );
  DFFQX1 dpl_reg_reg_2__6_ ( .D(N12590), .C(net12441), .Q(dpl_reg[22]) );
  DFFQX1 dpl_reg_reg_2__1_ ( .D(N12585), .C(net12441), .Q(dpl_reg[17]) );
  DFFQX1 dpl_reg_reg_2__0_ ( .D(N12584), .C(net12441), .Q(dpl_reg[16]) );
  DFFQX1 dph_reg_reg_6__7_ ( .D(N12555), .C(net12421), .Q(dph_reg[55]) );
  DFFQX1 dph_reg_reg_6__3_ ( .D(N12551), .C(net12421), .Q(dph_reg[51]) );
  DFFQX1 dph_reg_reg_6__1_ ( .D(N12549), .C(net12421), .Q(dph_reg[49]) );
  DFFQX1 dpl_reg_reg_6__7_ ( .D(N12627), .C(net12421), .Q(dpl_reg[55]) );
  DFFQX1 dpl_reg_reg_6__6_ ( .D(N12626), .C(net12421), .Q(dpl_reg[54]) );
  DFFQX1 dpl_reg_reg_6__1_ ( .D(N12621), .C(net12421), .Q(dpl_reg[49]) );
  DFFQX1 dpl_reg_reg_6__0_ ( .D(N12620), .C(net12421), .Q(dpl_reg[48]) );
  DFFQX1 ckcon_r_reg_3_ ( .D(N12968), .C(net12400), .Q(ckcon[3]) );
  DFFQX1 dec_accop_reg_17_ ( .D(N10580), .C(net12400), .Q(dec_accop[17]) );
  DFFQX1 ramwe_r_reg ( .D(N11487), .C(net12400), .Q(ramwe) );
  DFFQX1 pmw_reg_reg ( .D(n1939), .C(net12400), .Q(pmw) );
  DFFQX1 temp_reg_3_ ( .D(N12717), .C(net12496), .Q(temp[3]) );
  DFFQX1 temp_reg_4_ ( .D(N12718), .C(net12496), .Q(temp[4]) );
  DFFQX1 temp_reg_5_ ( .D(N12719), .C(net12496), .Q(temp[5]) );
  DFFQX1 temp_reg_6_ ( .D(N12720), .C(net12496), .Q(temp[6]) );
  DFFQX1 temp_reg_0_ ( .D(N12714), .C(net12496), .Q(temp[0]) );
  DFFQX1 temp_reg_1_ ( .D(N12715), .C(net12496), .Q(temp[1]) );
  DFFQX1 temp_reg_2_ ( .D(N12716), .C(net12496), .Q(temp[2]) );
  DFFQX1 temp_reg_7_ ( .D(N12721), .C(net12496), .Q(temp[7]) );
  DFFQX1 bitno_reg_0_ ( .D(N11492), .C(net12411), .Q(N343) );
  DFFQX1 bitno_reg_1_ ( .D(N11493), .C(net12411), .Q(N344) );
  DFFQX1 phase_reg_2_ ( .D(N681), .C(net12400), .Q(phase[2]) );
  DFFQX1 temp2_reg_6_ ( .D(N12729), .C(net12400), .Q(temp2_comb[6]) );
  DFFQX1 pc_reg_6_ ( .D(N486), .C(net12400), .Q(memaddr[6]) );
  DFFQX1 rn_reg_reg_19__3_ ( .D(n415), .C(net12601), .Q(rn_reg[99]) );
  DFFQX1 rn_reg_reg_27__3_ ( .D(n416), .C(net12641), .Q(rn_reg[35]) );
  DFFQX1 rn_reg_reg_16__3_ ( .D(n414), .C(net12586), .Q(rn_reg[123]) );
  DFFQX1 rn_reg_reg_20__3_ ( .D(n415), .C(net12606), .Q(rn_reg[91]) );
  DFFQX1 rn_reg_reg_24__3_ ( .D(n416), .C(net12626), .Q(rn_reg[59]) );
  DFFQX1 rn_reg_reg_28__3_ ( .D(n416), .C(net12646), .Q(rn_reg[27]) );
  DFFQX1 rn_reg_reg_17__3_ ( .D(n415), .C(net12591), .Q(rn_reg[115]) );
  DFFQX1 rn_reg_reg_21__3_ ( .D(n415), .C(net12611), .Q(rn_reg[83]) );
  DFFQX1 rn_reg_reg_25__3_ ( .D(n416), .C(net12631), .Q(rn_reg[51]) );
  DFFQX1 rn_reg_reg_29__3_ ( .D(n416), .C(net12651), .Q(rn_reg[19]) );
  DFFQX1 rn_reg_reg_18__3_ ( .D(n415), .C(net12596), .Q(rn_reg[107]) );
  DFFQX1 rn_reg_reg_26__3_ ( .D(n416), .C(net12636), .Q(rn_reg[43]) );
  DFFQX1 dps_reg_reg_2_ ( .D(N12695), .C(net12400), .Q(dps[2]) );
  DFFQX1 dec_accop_reg_11_ ( .D(N10574), .C(net12400), .Q(dec_accop[11]) );
  DFFQX1 dec_accop_reg_14_ ( .D(N10577), .C(net12400), .Q(dec_accop[14]) );
  DFFQX1 sp_reg_reg_0_ ( .D(N12697), .C(net12400), .Q(sp[0]) );
  DFFQX1 sp_reg_reg_1_ ( .D(N12698), .C(net12400), .Q(sp[1]) );
  DFFQX1 dec_accop_reg_12_ ( .D(N10575), .C(net12400), .Q(dec_accop[12]) );
  DFFQX1 dec_accop_reg_4_ ( .D(N10567), .C(net12400), .Q(dec_accop[4]) );
  DFFQX1 dec_accop_reg_3_ ( .D(N10566), .C(net12400), .Q(dec_accop[3]) );
  DFFQX1 rs_reg_reg_1_ ( .D(N12710), .C(net12400), .Q(rs[1]) );
  DFFQX1 dec_accop_reg_15_ ( .D(N10578), .C(net12400), .Q(dec_accop[15]) );
  DFFQX1 sp_reg_reg_2_ ( .D(N12699), .C(net12400), .Q(sp[2]) );
  DFFQX1 sfroe_r_reg ( .D(N11488), .C(net12400), .Q(sfroe_r) );
  DFFQX1 sfrwe_r_reg ( .D(N11489), .C(net12400), .Q(sfrwe_r) );
  DFFQX1 interrupt_reg ( .D(n1972), .C(net12406), .Q(interrupt) );
  DFFQX1 temp2_reg_5_ ( .D(N12728), .C(net12400), .Q(temp2_comb[5]) );
  DFFQX1 ramdatao_r_reg_4_ ( .D(N11502), .C(net12400), .Q(ramdatao[4]) );
  DFFQX1 ramdatao_r_reg_2_ ( .D(N11500), .C(net12400), .Q(ramdatao[2]) );
  DFFQX1 phase_reg_0_ ( .D(N679), .C(net12400), .Q(phase[0]) );
  DFFQX1 pc_reg_5_ ( .D(N485), .C(net12400), .Q(n2186) );
  DFFQX1 dec_accop_reg_13_ ( .D(N10576), .C(net12400), .Q(dec_accop[13]) );
  DFFQX1 dec_accop_reg_1_ ( .D(N10564), .C(net12400), .Q(dec_accop[1]) );
  DFFQX1 dec_accop_reg_0_ ( .D(N10563), .C(net12400), .Q(dec_accop[0]) );
  DFFQX1 dec_accop_reg_2_ ( .D(N10565), .C(net12400), .Q(dec_accop[2]) );
  DFFQX1 memrd_s_reg ( .D(N584), .C(net12400), .Q(memrd) );
  DFFQX1 accactv_reg ( .D(N10562), .C(net12400), .Q(accactv) );
  DFFQX1 waitcnt_reg_0_ ( .D(N12974), .C(net12501), .Q(waitcnt[0]) );
  DFFQX1 waitcnt_reg_1_ ( .D(N12975), .C(net12501), .Q(waitcnt[1]) );
  DFFQX1 ckcon_r_reg_0_ ( .D(N12965), .C(net12400), .Q(ckcon[0]) );
  DFFQX1 ckcon_r_reg_4_ ( .D(N12969), .C(net12400), .Q(ckcon[4]) );
  DFFQX1 ckcon_r_reg_5_ ( .D(N12970), .C(net12400), .Q(ckcon[5]) );
  DFFQX1 ckcon_r_reg_1_ ( .D(N12966), .C(net12400), .Q(ckcon[1]) );
  DFFQX1 ckcon_r_reg_2_ ( .D(N12967), .C(net12400), .Q(ckcon[2]) );
  DFFQX1 mempsrd_r_reg ( .D(N582), .C(net12400), .Q(mempsrd) );
  DFFQX1 mempswr_s_reg ( .D(N583), .C(net12400), .Q(mempswr) );
  DFFQX1 temp2_reg_4_ ( .D(N12727), .C(net12400), .Q(temp2_comb[4]) );
  DFFQX1 memwr_s_reg ( .D(N585), .C(net12400), .Q(memwr) );
  DFFQX1 acc_reg_reg_5_ ( .D(N12474), .C(net12400), .Q(acc[5]) );
  DFFQX1 acc_reg_reg_4_ ( .D(N12473), .C(net12400), .Q(acc[4]) );
  DFFQX1 instr_reg_2_ ( .D(N672), .C(net12406), .Q(n2193) );
  DFFQX1 pc_reg_15_ ( .D(N495), .C(net12400), .Q(pc_o[15]) );
  DFFQX1 phase_reg_1_ ( .D(N680), .C(net12400), .Q(phase[1]) );
  DFFQX1 acc_reg_reg_6_ ( .D(N12475), .C(net12400), .Q(acc[6]) );
  DFFQX1 pc_reg_14_ ( .D(N494), .C(net12400), .Q(memaddr[14]) );
  DFFQX1 pc_reg_3_ ( .D(N483), .C(net12400), .Q(pc_o[3]) );
  DFFQX1 pc_reg_4_ ( .D(N484), .C(net12400), .Q(n2187) );
  DFFQX1 instr_reg_4_ ( .D(N674), .C(net12406), .Q(n2191) );
  DFFQX1 instr_reg_0_ ( .D(N670), .C(net12406), .Q(N352) );
  DFFQX1 dps_reg_reg_1_ ( .D(N12694), .C(net12400), .Q(N350) );
  DFFQX1 dps_reg_reg_0_ ( .D(N12693), .C(net12400), .Q(dps[0]) );
  DFFQX1 rs_reg_reg_0_ ( .D(N12709), .C(net12400), .Q(rs[0]) );
  DFFQX1 dps_reg_reg_3_ ( .D(n1884), .C(net12400), .Q(dps[3]) );
  DFFQX1 waitcnt_reg_2_ ( .D(N12976), .C(net12501), .Q(waitcnt[2]) );
  DFFQX1 ckcon_r_reg_6_ ( .D(N12971), .C(net12400), .Q(ckcon[6]) );
  DFFQX1 temp2_reg_3_ ( .D(N12726), .C(net12400), .Q(temp2_comb[3]) );
  DFFQX1 instr_reg_7_ ( .D(N677), .C(net12406), .Q(n2188) );
  DFFQX1 ramdatao_r_reg_0_ ( .D(N11498), .C(net12400), .Q(ramdatao[0]) );
  DFFQX1 ramdatao_r_reg_1_ ( .D(N11499), .C(net12400), .Q(ramdatao[1]) );
  DFFQX1 instr_reg_1_ ( .D(N671), .C(net12406), .Q(n2194) );
  DFFQX1 pc_reg_11_ ( .D(N491), .C(net12400), .Q(pc_o[11]) );
  DFFQX1 pc_reg_12_ ( .D(N492), .C(net12400), .Q(memaddr[12]) );
  DFFQX1 pc_reg_2_ ( .D(N482), .C(net12400), .Q(pc_o[2]) );
  DFFQX1 pc_reg_8_ ( .D(N488), .C(net12400), .Q(memaddr[8]) );
  DFFQX1 pc_reg_10_ ( .D(N490), .C(net12400), .Q(pc_o[10]) );
  DFFQX1 pc_reg_9_ ( .D(N489), .C(net12400), .Q(pc_o[9]) );
  DFFQX1 instr_reg_3_ ( .D(N673), .C(net12406), .Q(n2192) );
  DFFQX1 pc_reg_13_ ( .D(N493), .C(net12400), .Q(pc_o[13]) );
  DFFQX1 pc_reg_7_ ( .D(N487), .C(net12400), .Q(n2185) );
  DFFQX1 ramsfrwe_reg ( .D(n1891), .C(net12400), .Q(ramsfrwe) );
  DFFQX1 instr_reg_5_ ( .D(N675), .C(net12406), .Q(n2190) );
  DFFQX1 ramsfraddr_s_reg_3_ ( .D(N11481), .C(net12400), .Q(ramsfraddr[3]) );
  DFFQX1 temp2_reg_1_ ( .D(N12724), .C(net12400), .Q(temp2_comb[1]) );
  DFFQX1 temp2_reg_2_ ( .D(N12725), .C(net12400), .Q(temp2_comb[2]) );
  DFFQX1 ramdatao_r_reg_3_ ( .D(N11501), .C(net12400), .Q(ramdatao[3]) );
  DFFQX1 instr_reg_6_ ( .D(N676), .C(net12406), .Q(n2189) );
  DFFQX1 pc_reg_0_ ( .D(N480), .C(net12400), .Q(N1761) );
  DFFQX1 pc_reg_1_ ( .D(N481), .C(net12400), .Q(pc_o[1]) );
  DFFQX1 divtempreg_reg_6_ ( .D(N13373), .C(net12671), .Q(divtempreg[6]) );
  DFFQX1 ac_reg_reg ( .D(N12706), .C(net12400), .Q(ac) );
  DFFQX1 divtempreg_reg_5_ ( .D(N13372), .C(net12671), .Q(divtempreg[5]) );
  DFFQX1 ramsfraddr_s_reg_1_ ( .D(N11479), .C(net12400), .Q(ramsfraddr[1]) );
  DFFQX1 ramsfraddr_s_reg_6_ ( .D(N11484), .C(net12400), .Q(ramsfraddr[6]) );
  DFFQX1 b_reg_reg_7_ ( .D(N12484), .C(net12400), .Q(b[7]) );
  DFFQX1 ramsfraddr_s_reg_2_ ( .D(N11480), .C(net12400), .Q(ramsfraddr[2]) );
  DFFQX1 ramsfraddr_s_reg_7_ ( .D(N11485), .C(net12400), .Q(ramsfraddr[7]) );
  DFFQX1 ramsfraddr_s_reg_0_ ( .D(N11478), .C(net12400), .Q(ramsfraddr[0]) );
  DFFQX1 ramsfraddr_s_reg_5_ ( .D(N11483), .C(net12400), .Q(ramsfraddr[5]) );
  DFFQX1 acc_reg_reg_3_ ( .D(N12472), .C(net12400), .Q(acc[3]) );
  DFFQX1 temp2_reg_0_ ( .D(N12723), .C(net12400), .Q(temp2_comb[0]) );
  DFFQX1 ramsfraddr_s_reg_4_ ( .D(N11482), .C(net12400), .Q(ramsfraddr[4]) );
  DFFQX1 acc_reg_reg_0_ ( .D(N12469), .C(net12400), .Q(acc[0]) );
  DFFQX1 dec_accop_reg_7_ ( .D(N10570), .C(net12400), .Q(dec_accop[7]) );
  DFFQX1 dec_accop_reg_8_ ( .D(N10571), .C(net12400), .Q(dec_accop[8]) );
  DFFQX1 dec_accop_reg_6_ ( .D(N10569), .C(net12400), .Q(dec_accop[6]) );
  DFFQX1 dec_accop_reg_16_ ( .D(N10579), .C(net12400), .Q(dec_accop[16]) );
  DFFQX1 dec_accop_reg_18_ ( .D(N10581), .C(net12400), .Q(dec_accop[18]) );
  DFFQX1 dec_accop_reg_9_ ( .D(N10572), .C(net12400), .Q(dec_accop[9]) );
  DFFQX1 divtempreg_reg_4_ ( .D(N13371), .C(net12671), .Q(divtempreg[4]) );
  DFFQX1 dec_accop_reg_5_ ( .D(N10568), .C(net12400), .Q(dec_accop[5]) );
  DFFQX1 c_reg_reg ( .D(N12705), .C(net12400), .Q(c) );
  DFFQX1 b_reg_reg_5_ ( .D(N12482), .C(net12400), .Q(b[5]) );
  DFFQX1 b_reg_reg_6_ ( .D(N12483), .C(net12400), .Q(b[6]) );
  DFFQX1 acc_reg_reg_2_ ( .D(N12471), .C(net12400), .Q(acc[2]) );
  DFFQX1 acc_reg_reg_1_ ( .D(N12470), .C(net12400), .Q(acc[1]) );
  DFFQX1 divtempreg_reg_2_ ( .D(N13369), .C(net12671), .Q(divtempreg[2]) );
  DFFQX1 divtempreg_reg_3_ ( .D(N13370), .C(net12671), .Q(divtempreg[3]) );
  DFFQX1 dec_accop_reg_10_ ( .D(N10573), .C(net12400), .Q(dec_accop[10]) );
  DFFQX1 b_reg_reg_4_ ( .D(N12481), .C(net12400), .Q(b[4]) );
  DFFQX1 divtempreg_reg_1_ ( .D(N13368), .C(net12671), .Q(divtempreg[1]) );
  DFFQX1 b_reg_reg_3_ ( .D(N12480), .C(net12400), .Q(b[3]) );
  DFFQX1 divtempreg_reg_0_ ( .D(N13367), .C(net12671), .Q(divtempreg[0]) );
  DFFQX1 b_reg_reg_1_ ( .D(N12478), .C(net12400), .Q(b[1]) );
  DFFQX1 b_reg_reg_0_ ( .D(N12477), .C(net12400), .Q(b[0]) );
  DFFQX1 acc_reg_reg_7_ ( .D(N12476), .C(net12400), .Q(acc[7]) );
  DFFQX1 b_reg_reg_2_ ( .D(N12479), .C(net12400), .Q(b[2]) );
  INVXL U3 ( .A(n1554), .Y(n1561) );
  OAI222X1 U4 ( .A(n676), .B(n1352), .C(n871), .D(n675), .E(n2173), .F(n674), 
        .Y(n741) );
  OAI222X1 U5 ( .A(n676), .B(n1564), .C(n1566), .D(n675), .E(n2167), .F(n674), 
        .Y(n1574) );
  NOR2X2 U6 ( .A(n1475), .B(n382), .Y(n146) );
  NOR21XL U7 ( .B(cpu_hold), .A(n1940), .Y(n735) );
  INVX2 U8 ( .A(n1272), .Y(n1065) );
  NAND3X1 U9 ( .A(n136), .B(n137), .C(n138), .Y(n1302) );
  NAND3X1 U10 ( .A(n133), .B(n134), .C(n135), .Y(n1404) );
  NAND21X1 U11 ( .B(n430), .A(n572), .Y(n573) );
  NAND3X1 U12 ( .A(n130), .B(n131), .C(n132), .Y(n1419) );
  AO21X1 U13 ( .B(n542), .C(n1365), .A(n1225), .Y(n543) );
  INVX1 U14 ( .A(sfrdatai[6]), .Y(n1547) );
  INVX1 U15 ( .A(sfrdatai[5]), .Y(n1544) );
  INVX1 U16 ( .A(n1292), .Y(n766) );
  MUX2X1 U17 ( .D0(memaddr[6]), .D1(n1484), .S(n146), .Y(memaddr_comb[6]) );
  OR2X1 U18 ( .A(n2087), .B(n916), .Y(n4) );
  AO21X1 U19 ( .B(n2118), .C(n2036), .A(n1480), .Y(n5) );
  OA222X1 U20 ( .A(n1352), .B(n1563), .C(n871), .D(n1565), .E(n2173), .F(n192), 
        .Y(n6) );
  OA21X1 U21 ( .B(n1810), .C(n1809), .A(n1811), .Y(n7) );
  OR4X1 U22 ( .A(n2131), .B(ramsfraddr[5]), .C(ramsfraddr[6]), .D(
        ramsfraddr[7]), .Y(n8) );
  INVXL U23 ( .A(n1682), .Y(n9) );
  INVXL U24 ( .A(n9), .Y(n10) );
  INVXL U28 ( .A(n804), .Y(n11) );
  INVXL U29 ( .A(n804), .Y(n12) );
  INVXL U30 ( .A(n805), .Y(n13) );
  INVXL U31 ( .A(n805), .Y(n14) );
  INVXL U32 ( .A(n2089), .Y(n15) );
  INVXL U33 ( .A(n15), .Y(n16) );
  INVXL U34 ( .A(pc_o[15]), .Y(n17) );
  INVXL U35 ( .A(n17), .Y(memaddr[15]) );
  INVXL U36 ( .A(n2189), .Y(n19) );
  INVXL U37 ( .A(n19), .Y(instr[6]) );
  INVXL U38 ( .A(n1499), .Y(n21) );
  INVXL U39 ( .A(n1499), .Y(n22) );
  INVXL U40 ( .A(n2186), .Y(n23) );
  INVXL U41 ( .A(n23), .Y(pc_o[5]) );
  INVXL U42 ( .A(memaddr[6]), .Y(n25) );
  INVXL U43 ( .A(n25), .Y(pc_o[6]) );
  INVXL U44 ( .A(pc_o[10]), .Y(n27) );
  INVXL U45 ( .A(n27), .Y(memaddr[10]) );
  INVXL U46 ( .A(pc_o[11]), .Y(n29) );
  INVXL U47 ( .A(n29), .Y(memaddr[11]) );
  INVXL U48 ( .A(memaddr[8]), .Y(n31) );
  INVXL U49 ( .A(n31), .Y(pc_o[8]) );
  INVXL U50 ( .A(pc_o[2]), .Y(n33) );
  INVXL U51 ( .A(n33), .Y(memaddr[2]) );
  INVXL U52 ( .A(memaddr[12]), .Y(n35) );
  INVXL U53 ( .A(n35), .Y(pc_o[12]) );
  INVXL U54 ( .A(N1761), .Y(n37) );
  INVXL U55 ( .A(n37), .Y(memaddr[0]) );
  INVXL U56 ( .A(pc_o[9]), .Y(n39) );
  INVXL U57 ( .A(n39), .Y(memaddr[9]) );
  INVXL U58 ( .A(memaddr[14]), .Y(n41) );
  INVXL U59 ( .A(n41), .Y(pc_o[14]) );
  INVXL U60 ( .A(pc_o[1]), .Y(n43) );
  INVXL U61 ( .A(n43), .Y(memaddr[1]) );
  INVXL U62 ( .A(pc_o[3]), .Y(n45) );
  INVXL U63 ( .A(n45), .Y(memaddr[3]) );
  INVXL U64 ( .A(pc_o[13]), .Y(n47) );
  INVXL U65 ( .A(n47), .Y(memaddr[13]) );
  INVXL U66 ( .A(n47), .Y(n49) );
  INVXL U67 ( .A(n2185), .Y(n50) );
  INVXL U68 ( .A(n50), .Y(memaddr[7]) );
  INVXL U69 ( .A(n50), .Y(pc_o[7]) );
  INVXL U70 ( .A(n2187), .Y(n53) );
  INVXL U71 ( .A(n53), .Y(memaddr[4]) );
  INVXL U72 ( .A(n53), .Y(pc_o[4]) );
  BUFX3 U73 ( .A(n2039), .Y(n56) );
  INVX1 U74 ( .A(instr[7]), .Y(n57) );
  BUFX3 U75 ( .A(n1258), .Y(n58) );
  BUFX3 U76 ( .A(n2188), .Y(instr[7]) );
  BUFX3 U77 ( .A(n1260), .Y(n60) );
  INVX1 U78 ( .A(n64), .Y(instr[2]) );
  BUFX3 U79 ( .A(n1262), .Y(n62) );
  BUFX3 U80 ( .A(n1955), .Y(n63) );
  BUFX3 U81 ( .A(n2106), .Y(n64) );
  BUFX3 U82 ( .A(n1267), .Y(n65) );
  BUFX3 U83 ( .A(n1250), .Y(n66) );
  AOI21X1 U84 ( .B(n1634), .C(n178), .A(n396), .Y(n1251) );
  INVX1 U85 ( .A(n1251), .Y(n67) );
  INVX1 U86 ( .A(n1251), .Y(n68) );
  INVX1 U87 ( .A(instr[1]), .Y(n69) );
  INVX1 U88 ( .A(n1966), .Y(n70) );
  BUFX3 U89 ( .A(n2194), .Y(instr[1]) );
  AOI21X1 U90 ( .B(n385), .C(n155), .A(n1808), .Y(n1257) );
  INVX1 U91 ( .A(n1257), .Y(n72) );
  INVX1 U92 ( .A(n1257), .Y(n73) );
  AOI21X1 U93 ( .B(n1634), .C(n180), .A(n398), .Y(n1249) );
  INVX1 U94 ( .A(n1249), .Y(n74) );
  INVX1 U95 ( .A(n1249), .Y(n75) );
  BUFX3 U96 ( .A(n1252), .Y(n76) );
  NOR2X1 U97 ( .A(n1329), .B(n1244), .Y(n1266) );
  INVX1 U98 ( .A(n1266), .Y(n77) );
  INVX1 U99 ( .A(n1266), .Y(n78) );
  INVX1 U100 ( .A(n810), .Y(n79) );
  INVX1 U101 ( .A(n2044), .Y(n80) );
  AOI21X1 U102 ( .B(n385), .C(n154), .A(n396), .Y(n1259) );
  INVX1 U103 ( .A(n1259), .Y(n81) );
  INVX1 U104 ( .A(n1259), .Y(n82) );
  BUFX3 U105 ( .A(n1254), .Y(n83) );
  AOI21X1 U106 ( .B(n1634), .C(n181), .A(n396), .Y(n1255) );
  INVX1 U107 ( .A(n1255), .Y(n84) );
  INVX1 U108 ( .A(n1255), .Y(n85) );
  INVX1 U109 ( .A(n615), .Y(n86) );
  BUFX3 U110 ( .A(n1269), .Y(n87) );
  NAND2X1 U111 ( .A(n1015), .B(n1942), .Y(n88) );
  INVX1 U112 ( .A(n2192), .Y(n89) );
  INVX1 U113 ( .A(n815), .Y(n90) );
  NAND2X1 U114 ( .A(n1014), .B(n1942), .Y(n91) );
  INVX1 U115 ( .A(n519), .Y(n92) );
  AOI21X1 U116 ( .B(n385), .C(n152), .A(n398), .Y(n1263) );
  INVX1 U117 ( .A(n1263), .Y(n93) );
  INVX1 U118 ( .A(n1263), .Y(n94) );
  AOI21X1 U119 ( .B(n1634), .C(n179), .A(n397), .Y(n1253) );
  INVX1 U120 ( .A(n1253), .Y(n95) );
  INVX1 U121 ( .A(n1253), .Y(n96) );
  BUFX3 U122 ( .A(n1256), .Y(n97) );
  NOR2X1 U123 ( .A(n1326), .B(n1244), .Y(n98) );
  INVX1 U124 ( .A(n614), .Y(n99) );
  NAND2X1 U125 ( .A(n1747), .B(n2193), .Y(N354) );
  INVX1 U126 ( .A(N354), .Y(n100) );
  INVX1 U127 ( .A(N354), .Y(n101) );
  INVX1 U128 ( .A(n123), .Y(n102) );
  INVX1 U129 ( .A(n2192), .Y(n103) );
  INVX1 U130 ( .A(n103), .Y(n104) );
  INVX1 U131 ( .A(n103), .Y(instr[3]) );
  INVX1 U132 ( .A(n2127), .Y(n106) );
  BUFX3 U133 ( .A(n1709), .Y(n107) );
  AOI21X1 U134 ( .B(n385), .C(n153), .A(n398), .Y(n1261) );
  INVX1 U135 ( .A(n1261), .Y(n108) );
  INVX1 U136 ( .A(n1261), .Y(n109) );
  BUFX3 U137 ( .A(n1264), .Y(n110) );
  NOR2X1 U138 ( .A(n1325), .B(n1244), .Y(n111) );
  INVX1 U139 ( .A(n783), .Y(n112) );
  NAND2X1 U140 ( .A(n806), .B(n808), .Y(n113) );
  INVX1 U141 ( .A(n1189), .Y(n114) );
  MUX4X1 U142 ( .D0(n362), .D1(n360), .D2(n361), .D3(n359), .S0(n2065), .S1(
        n100), .Y(n363) );
  INVX1 U143 ( .A(accactv), .Y(n383) );
  INVX1 U144 ( .A(n383), .Y(n115) );
  INVX1 U145 ( .A(n383), .Y(n116) );
  INVX1 U146 ( .A(N348), .Y(n117) );
  INVX1 U147 ( .A(n117), .Y(n118) );
  INVX1 U148 ( .A(n117), .Y(n119) );
  OAI221X1 U149 ( .A(n1335), .B(n441), .C(n1188), .D(n1336), .E(n1341), .Y(
        N348) );
  INVX1 U150 ( .A(n2191), .Y(n120) );
  INVX1 U151 ( .A(n120), .Y(n121) );
  INVX1 U152 ( .A(n120), .Y(instr[4]) );
  BUFX3 U153 ( .A(phase[0]), .Y(n2103) );
  INVX1 U154 ( .A(n2103), .Y(n123) );
  INVX1 U155 ( .A(n2103), .Y(n124) );
  INVX1 U156 ( .A(n2103), .Y(n125) );
  INVX1 U157 ( .A(n382), .Y(waitstaten) );
  OR2X2 U158 ( .A(n676), .B(n965), .Y(n127) );
  OR2X1 U159 ( .A(n1131), .B(n675), .Y(n128) );
  OR2X1 U160 ( .A(n674), .B(n648), .Y(n129) );
  NAND3X1 U161 ( .A(n127), .B(n128), .C(n129), .Y(n669) );
  INVX3 U162 ( .A(n959), .Y(n1475) );
  NAND21X1 U163 ( .B(n1961), .A(n647), .Y(n676) );
  OR2X1 U164 ( .A(n676), .B(n1544), .Y(n130) );
  OR2X1 U165 ( .A(n847), .B(n675), .Y(n131) );
  OR2X1 U166 ( .A(n2169), .B(n674), .Y(n132) );
  NAND2XL U167 ( .A(n675), .B(n676), .Y(n674) );
  OR2X1 U168 ( .A(n676), .B(n1343), .Y(n136) );
  OR2X1 U169 ( .A(n2038), .B(n647), .Y(n675) );
  OR2X1 U170 ( .A(n676), .B(n1541), .Y(n133) );
  OR2X1 U171 ( .A(n853), .B(n675), .Y(n134) );
  OR2XL U172 ( .A(n2170), .B(n674), .Y(n135) );
  INVX1 U173 ( .A(sfrdatai[4]), .Y(n1541) );
  NAND42X1 U174 ( .C(n472), .D(n469), .A(n466), .B(n465), .Y(n1399) );
  NOR2X1 U175 ( .A(n1475), .B(n382), .Y(n145) );
  INVX1 U176 ( .A(sfrdatai[2]), .Y(n1343) );
  OR2X1 U177 ( .A(n2172), .B(n674), .Y(n138) );
  OR2X1 U178 ( .A(n865), .B(n675), .Y(n137) );
  INVXL U179 ( .A(n1302), .Y(n1322) );
  AO21XL U180 ( .B(n752), .C(n660), .A(n1523), .Y(n754) );
  INVXL U181 ( .A(n669), .Y(n665) );
  NAND21XL U182 ( .B(n1584), .A(n665), .Y(n649) );
  OAI222XL U183 ( .A(n676), .B(n1547), .C(n841), .D(n675), .E(n2168), .F(n674), 
        .Y(n1554) );
  AND2XL U184 ( .A(n400), .B(n1086), .Y(N12469) );
  AND2XL U185 ( .A(n390), .B(n983), .Y(N12470) );
  NOR32XL U186 ( .B(n1526), .C(n1421), .A(n139), .Y(n746) );
  MUX2IX1 U187 ( .D0(n1584), .D1(n1576), .S(n172), .Y(n139) );
  OAI222XL U188 ( .A(n965), .B(n1563), .C(n1131), .D(n1565), .E(n192), .F(n648), .Y(n755) );
  XNOR3X1 U189 ( .A(n140), .B(n1570), .C(n1569), .Y(incdec_out[7]) );
  OAI222XL U190 ( .A(n2167), .B(n192), .C(n1566), .D(n1565), .E(n1564), .F(
        n1563), .Y(n140) );
  NAND31XL U191 ( .C(n469), .A(memack), .B(n468), .Y(n1710) );
  INVX1 U192 ( .A(n735), .Y(n182) );
  MUX2AXL U193 ( .D0(n141), .D1(pdmode), .S(n1290), .Y(n1973) );
  OAI21X1 U194 ( .B(codefetch_s), .C(n1273), .A(n457), .Y(n141) );
  OAI31XL U195 ( .A(n768), .B(n2019), .C(n1840), .D(mempsrd), .Y(n1804) );
  OAI222XL U196 ( .A(n124), .B(n715), .C(n2078), .D(n716), .E(n1675), .F(n2077), .Y(n1297) );
  NOR3XL U197 ( .A(n2071), .B(ramsfraddr[2]), .C(n2119), .Y(n1015) );
  OR2X1 U198 ( .A(n676), .B(n1534), .Y(n142) );
  OR2X1 U199 ( .A(n1533), .B(n675), .Y(n143) );
  OR2X1 U200 ( .A(n2171), .B(n674), .Y(n144) );
  NAND3X1 U201 ( .A(n142), .B(n143), .C(n144), .Y(n1519) );
  INVX1 U202 ( .A(sfrdatai[3]), .Y(n1534) );
  INVX1 U203 ( .A(n397), .Y(n387) );
  INVX1 U204 ( .A(n397), .Y(n388) );
  INVX1 U205 ( .A(n398), .Y(n389) );
  INVX1 U206 ( .A(n396), .Y(n393) );
  INVX1 U207 ( .A(n396), .Y(n394) );
  INVX1 U208 ( .A(n1808), .Y(n395) );
  INVX1 U209 ( .A(n396), .Y(n391) );
  INVX1 U210 ( .A(n396), .Y(n390) );
  INVX1 U211 ( .A(n396), .Y(n392) );
  INVX1 U212 ( .A(n437), .Y(n285) );
  INVX1 U213 ( .A(n652), .Y(n654) );
  INVX1 U214 ( .A(n401), .Y(n397) );
  INVX1 U215 ( .A(n400), .Y(n398) );
  INVX1 U216 ( .A(n400), .Y(n396) );
  NAND21X1 U217 ( .B(n450), .A(n452), .Y(N370) );
  INVX1 U218 ( .A(n400), .Y(n399) );
  INVX1 U219 ( .A(n435), .Y(n287) );
  INVX1 U220 ( .A(n437), .Y(n286) );
  INVX1 U221 ( .A(n607), .Y(n545) );
  INVX1 U222 ( .A(n1575), .Y(n2038) );
  INVX1 U223 ( .A(n1409), .Y(n2045) );
  INVX1 U224 ( .A(n2036), .Y(n1908) );
  NAND21X1 U225 ( .B(n1573), .A(n1575), .Y(n652) );
  INVX1 U226 ( .A(n1521), .Y(n653) );
  INVX1 U227 ( .A(n2007), .Y(n425) );
  INVX1 U228 ( .A(n2006), .Y(n421) );
  INVX1 U229 ( .A(n2005), .Y(n417) );
  INVX1 U230 ( .A(n1808), .Y(n401) );
  INVX1 U231 ( .A(n2007), .Y(n428) );
  INVX1 U232 ( .A(n2006), .Y(n424) );
  INVX1 U233 ( .A(n2005), .Y(n420) );
  INVX1 U234 ( .A(n2000), .Y(n404) );
  INVX1 U235 ( .A(n2001), .Y(n407) );
  INVX1 U236 ( .A(n2004), .Y(n416) );
  INVX1 U237 ( .A(n2003), .Y(n413) );
  INVX1 U238 ( .A(n2007), .Y(n427) );
  INVX1 U239 ( .A(n2006), .Y(n423) );
  INVX1 U240 ( .A(n2005), .Y(n419) );
  INVX1 U241 ( .A(n2002), .Y(n410) );
  INVX1 U242 ( .A(n2000), .Y(n403) );
  INVX1 U243 ( .A(n2007), .Y(n426) );
  INVX1 U244 ( .A(n2006), .Y(n422) );
  INVX1 U245 ( .A(n2005), .Y(n418) );
  INVX1 U246 ( .A(n2004), .Y(n415) );
  INVX1 U247 ( .A(n2003), .Y(n412) );
  INVX1 U248 ( .A(n2002), .Y(n409) );
  INVX1 U249 ( .A(n2001), .Y(n406) );
  INVX1 U250 ( .A(n1808), .Y(n400) );
  AND2X1 U251 ( .A(n391), .B(n1453), .Y(N11482) );
  AND2X1 U252 ( .A(n392), .B(n1454), .Y(N11484) );
  INVX1 U253 ( .A(n459), .Y(n452) );
  INVX1 U254 ( .A(n458), .Y(n453) );
  INVX1 U255 ( .A(n459), .Y(n454) );
  INVX1 U256 ( .A(n458), .Y(n455) );
  INVX1 U257 ( .A(n458), .Y(n456) );
  INVX1 U258 ( .A(n458), .Y(n457) );
  NAND21X1 U259 ( .B(n1523), .A(n649), .Y(n650) );
  INVXL U260 ( .A(n741), .Y(n752) );
  INVX1 U261 ( .A(n1293), .Y(n981) );
  INVX1 U262 ( .A(n437), .Y(n436) );
  NAND21X1 U263 ( .B(n917), .A(n1947), .Y(n2034) );
  MUX2X1 U264 ( .D0(n1576), .D1(n1584), .S(n1561), .Y(n1558) );
  NOR2X1 U265 ( .A(n2047), .B(n2046), .Y(n1409) );
  INVX1 U266 ( .A(n435), .Y(n288) );
  INVX1 U267 ( .A(n524), .Y(n1920) );
  INVX1 U268 ( .A(n975), .Y(n956) );
  INVX1 U269 ( .A(n1519), .Y(n1524) );
  NAND3X1 U270 ( .A(n1363), .B(n1364), .C(n1951), .Y(n607) );
  NAND21X1 U271 ( .B(n430), .A(n1156), .Y(n1575) );
  MUX2X1 U272 ( .D0(n1576), .D1(n1584), .S(n1322), .Y(n1334) );
  INVX1 U273 ( .A(n2037), .Y(n1947) );
  INVX1 U274 ( .A(n438), .Y(n250) );
  INVX1 U275 ( .A(n438), .Y(n252) );
  INVX1 U276 ( .A(n440), .Y(n246) );
  INVX1 U277 ( .A(n440), .Y(n248) );
  INVX1 U278 ( .A(n488), .Y(n1927) );
  OAI21X1 U279 ( .B(n431), .C(n1726), .A(n658), .Y(n1730) );
  INVX1 U280 ( .A(n438), .Y(n249) );
  INVX1 U281 ( .A(n1971), .Y(n1886) );
  INVX1 U282 ( .A(n917), .Y(n1952) );
  NOR2X1 U283 ( .A(n1995), .B(n727), .Y(N673) );
  NOR2X1 U284 ( .A(n1996), .B(n727), .Y(N674) );
  NOR2X1 U285 ( .A(n1998), .B(n727), .Y(N676) );
  INVX1 U286 ( .A(n1200), .Y(n1951) );
  NAND3X1 U287 ( .A(n666), .B(n690), .C(n573), .Y(n2036) );
  INVX1 U288 ( .A(n438), .Y(n251) );
  INVX1 U289 ( .A(n608), .Y(n2048) );
  INVX1 U290 ( .A(n441), .Y(n245) );
  INVX1 U291 ( .A(n441), .Y(n244) );
  INVX1 U292 ( .A(n628), .Y(n623) );
  INVX1 U293 ( .A(n440), .Y(n247) );
  INVX1 U294 ( .A(n577), .Y(n992) );
  NAND21X1 U295 ( .B(n2042), .A(n1911), .Y(n577) );
  INVX1 U296 ( .A(n574), .Y(n1021) );
  NAND21X1 U297 ( .B(n575), .A(n442), .Y(n574) );
  INVX1 U298 ( .A(n1196), .Y(n769) );
  INVX1 U299 ( .A(n625), .Y(n630) );
  NAND21X1 U300 ( .B(n624), .A(n623), .Y(n625) );
  INVX1 U301 ( .A(n719), .Y(n1016) );
  NAND21X1 U302 ( .B(n978), .A(n4), .Y(n719) );
  INVX1 U303 ( .A(n2087), .Y(n1946) );
  INVX1 U304 ( .A(n614), .Y(n620) );
  NAND32X1 U305 ( .B(n575), .C(n369), .A(n1907), .Y(n1585) );
  NAND32X1 U306 ( .B(n579), .C(n652), .A(n1572), .Y(n1480) );
  INVX1 U307 ( .A(n668), .Y(n579) );
  INVX1 U308 ( .A(n590), .Y(n1356) );
  NAND3X1 U309 ( .A(n2034), .B(n1600), .C(n1601), .Y(n1573) );
  NAND2X1 U310 ( .A(n2041), .B(n1061), .Y(n1601) );
  INVX1 U311 ( .A(n909), .Y(n505) );
  NAND21X1 U312 ( .B(n655), .A(n654), .Y(n1576) );
  NAND32X1 U313 ( .B(n1573), .C(n1156), .A(n1008), .Y(n923) );
  NAND21X1 U314 ( .B(n1909), .A(n644), .Y(n707) );
  INVX1 U315 ( .A(n1458), .Y(n1905) );
  INVX1 U316 ( .A(n569), .Y(n1008) );
  NAND21X1 U317 ( .B(n782), .A(n717), .Y(n569) );
  NOR2X1 U318 ( .A(n2094), .B(n2087), .Y(n977) );
  INVX1 U319 ( .A(n921), .Y(n781) );
  INVX1 U320 ( .A(n1686), .Y(n2094) );
  INVX1 U321 ( .A(n1640), .Y(n2091) );
  NAND21X1 U322 ( .B(n1904), .A(n450), .Y(n1450) );
  OR2X1 U323 ( .A(n652), .B(n651), .Y(n1521) );
  INVX1 U324 ( .A(n1456), .Y(n1909) );
  INVX1 U325 ( .A(n1572), .Y(n1523) );
  INVX1 U326 ( .A(n386), .Y(n384) );
  INVX1 U327 ( .A(n386), .Y(n385) );
  INVX1 U328 ( .A(n809), .Y(n1945) );
  INVX1 U329 ( .A(n885), .Y(n1027) );
  NAND21X1 U330 ( .B(rst), .A(waitstaten), .Y(n1808) );
  INVX1 U331 ( .A(n2002), .Y(n408) );
  INVX1 U332 ( .A(n2001), .Y(n405) );
  INVX1 U333 ( .A(n2003), .Y(n411) );
  INVX1 U334 ( .A(n2004), .Y(n414) );
  INVX1 U335 ( .A(n662), .Y(n1453) );
  NAND21X1 U336 ( .B(n1641), .A(n152), .Y(n1264) );
  NAND21X1 U337 ( .B(n1641), .A(n153), .Y(n1262) );
  NAND21X1 U338 ( .B(n1641), .A(n154), .Y(n1260) );
  NAND21X1 U339 ( .B(n1641), .A(n155), .Y(n1258) );
  NAND21X1 U340 ( .B(n386), .A(n387), .Y(n1641) );
  INVX1 U341 ( .A(n1020), .Y(N11494) );
  NAND21X1 U342 ( .B(n1993), .A(n389), .Y(n1020) );
  INVX1 U343 ( .A(n613), .Y(n616) );
  NAND21X1 U344 ( .B(n1307), .A(n614), .Y(n613) );
  AO21X1 U345 ( .B(n395), .C(n155), .A(n461), .Y(N12520) );
  AO21X1 U346 ( .B(n395), .C(n154), .A(n461), .Y(N12511) );
  AO21X1 U347 ( .B(n400), .C(n153), .A(n461), .Y(N12502) );
  AO21X1 U348 ( .B(n400), .C(n152), .A(n461), .Y(N12493) );
  INVX1 U349 ( .A(n661), .Y(n1454) );
  INVX1 U350 ( .A(n2000), .Y(n402) );
  INVX1 U351 ( .A(n811), .Y(n743) );
  INVX1 U352 ( .A(n1019), .Y(N11493) );
  NAND21X1 U353 ( .B(n1992), .A(n389), .Y(n1019) );
  INVX1 U354 ( .A(n1033), .Y(N10580) );
  NAND21X1 U355 ( .B(n1764), .A(n389), .Y(n1033) );
  INVX1 U356 ( .A(n1018), .Y(N11492) );
  NAND21X1 U357 ( .B(n1991), .A(n389), .Y(n1018) );
  OA21X1 U358 ( .B(n1027), .C(n150), .A(n394), .Y(N10572) );
  AND2X1 U359 ( .A(n1711), .B(n393), .Y(N11483) );
  AND2X1 U360 ( .A(n391), .B(n1452), .Y(N11481) );
  NOR21XL U361 ( .B(n390), .A(n1761), .Y(N10583) );
  NOR21XL U362 ( .B(n390), .A(n1762), .Y(N10582) );
  NOR21XL U363 ( .B(n400), .A(n1756), .Y(N10589) );
  NOR21XL U364 ( .B(n390), .A(n1805), .Y(N10564) );
  NOR21XL U365 ( .B(n400), .A(n1802), .Y(N10567) );
  NOR21XL U366 ( .B(n401), .A(n1767), .Y(N10577) );
  NOR21XL U367 ( .B(n401), .A(n1801), .Y(N10568) );
  AND2X1 U368 ( .A(n1887), .B(n393), .Y(N10588) );
  AND2X1 U369 ( .A(n1890), .B(n392), .Y(N10565) );
  NOR21XL U370 ( .B(n390), .A(n1806), .Y(N10563) );
  NOR21XL U371 ( .B(n390), .A(n1166), .Y(N10585) );
  INVX1 U372 ( .A(n818), .Y(n1198) );
  AOI31X1 U373 ( .A(n716), .B(n1016), .C(n1008), .D(n399), .Y(N690) );
  INVX1 U374 ( .A(n997), .Y(n1891) );
  INVX1 U375 ( .A(n1468), .Y(n2079) );
  NOR3XL U376 ( .A(n1072), .B(n22), .C(n1071), .Y(n1103) );
  INVX1 U377 ( .A(n1068), .Y(n2026) );
  NOR31X1 U378 ( .C(n1756), .A(n1784), .B(n1785), .Y(n1837) );
  AND2X1 U379 ( .A(n1737), .B(n1922), .Y(n1796) );
  AND2X1 U380 ( .A(n1061), .B(n1686), .Y(n1784) );
  INVX1 U381 ( .A(n1094), .Y(n2024) );
  NAND2X1 U382 ( .A(n2070), .B(n452), .Y(n1030) );
  INVX1 U383 ( .A(n463), .Y(n458) );
  INVX1 U384 ( .A(n463), .Y(n459) );
  NOR2X1 U385 ( .A(n458), .B(n2067), .Y(n687) );
  INVX1 U386 ( .A(n457), .Y(n461) );
  INVX1 U387 ( .A(n457), .Y(n460) );
  INVX1 U388 ( .A(n457), .Y(n462) );
  MUX2BXL U389 ( .D0(memwr), .D1(n1459), .S(waitstaten), .Y(memwr_comb) );
  NAND2X1 U390 ( .A(n755), .B(n756), .Y(n1353) );
  OR2X1 U391 ( .A(n1537), .B(n147), .Y(n706) );
  XNOR2XL U392 ( .A(n755), .B(n756), .Y(n147) );
  INVX1 U393 ( .A(n1399), .Y(n2184) );
  NOR2XL U394 ( .A(n1475), .B(n974), .Y(n148) );
  NOR2XL U395 ( .A(n1475), .B(n973), .Y(n149) );
  NAND21X1 U396 ( .B(n846), .A(n823), .Y(n1161) );
  OAI222XL U397 ( .A(n1700), .B(n1995), .C(n1701), .D(n724), .E(n1712), .F(
        n1998), .Y(n1452) );
  INVX1 U398 ( .A(n1041), .Y(n724) );
  OAI221X1 U399 ( .A(n1038), .B(n1701), .C(n1700), .D(n1997), .E(n1712), .Y(
        n1711) );
  NAND5XL U400 ( .A(n662), .B(n661), .C(sfrwe_comb_s), .D(n732), .E(n731), .Y(
        n1293) );
  INVX1 U401 ( .A(n1452), .Y(n732) );
  AND4X1 U402 ( .A(n1451), .B(n157), .C(n156), .D(n729), .Y(n731) );
  INVX1 U403 ( .A(n1711), .Y(n729) );
  GEN2XL U404 ( .D(n779), .E(n777), .C(n776), .B(n774), .A(n773), .Y(n803) );
  INVX1 U405 ( .A(n796), .Y(n774) );
  INVX1 U406 ( .A(n949), .Y(n773) );
  MUX2X1 U407 ( .D0(n1911), .D1(n772), .S(n158), .Y(n776) );
  NAND21X1 U408 ( .B(n79), .A(n844), .Y(n838) );
  INVX1 U409 ( .A(n816), .Y(n821) );
  NAND32X1 U410 ( .B(n838), .C(n818), .A(n815), .Y(n816) );
  INVX1 U411 ( .A(n814), .Y(n844) );
  NAND21X1 U412 ( .B(n1160), .A(n386), .Y(n814) );
  INVX1 U413 ( .A(memdatai[7]), .Y(n1999) );
  INVX1 U414 ( .A(n1455), .Y(n1298) );
  OA22X1 U415 ( .A(n1700), .B(n1998), .C(n1042), .D(n1701), .Y(n661) );
  AOI22BXL U416 ( .B(n1700), .A(memdatai[4]), .D(n1701), .C(n1045), .Y(n662)
         );
  INVX1 U417 ( .A(memdatai[1]), .Y(n1992) );
  INVX1 U418 ( .A(memdatai[3]), .Y(n1995) );
  INVX1 U419 ( .A(memdatai[6]), .Y(n1998) );
  INVX1 U420 ( .A(memdatai[4]), .Y(n1996) );
  INVX1 U421 ( .A(memdatai[5]), .Y(n1997) );
  INVX1 U422 ( .A(memdatai[0]), .Y(n1991) );
  INVX1 U423 ( .A(memdatai[2]), .Y(n1993) );
  XNOR2XL U424 ( .A(n1230), .B(n2062), .Y(n1231) );
  AOI22BXL U425 ( .B(n1230), .A(N11560), .D(n1231), .C(n1232), .Y(n1184) );
  INVX1 U426 ( .A(n1075), .Y(n1885) );
  INVX1 U427 ( .A(N11560), .Y(n2062) );
  INVX1 U428 ( .A(n1381), .Y(n2114) );
  NAND2X1 U429 ( .A(n843), .B(n844), .Y(n975) );
  NAND21X1 U430 ( .B(n846), .A(n845), .Y(n976) );
  INVX1 U431 ( .A(n839), .Y(n845) );
  NAND32X1 U432 ( .B(n838), .C(n843), .A(n837), .Y(n839) );
  INVX1 U433 ( .A(n435), .Y(n434) );
  INVX1 U434 ( .A(n877), .Y(n971) );
  INVX1 U435 ( .A(N346), .Y(n437) );
  INVX1 U436 ( .A(n1340), .Y(n2074) );
  INVX1 U437 ( .A(n1168), .Y(n2067) );
  INVX1 U438 ( .A(n1338), .Y(n2075) );
  INVX1 U439 ( .A(n1604), .Y(n1434) );
  INVX1 U440 ( .A(n1535), .Y(n1359) );
  XNOR2XL U441 ( .A(n1041), .B(n1045), .Y(n1046) );
  INVX1 U442 ( .A(n375), .Y(n379) );
  INVX1 U443 ( .A(n375), .Y(n378) );
  AOI33X1 U444 ( .A(n1038), .B(n1990), .C(n1039), .D(n1040), .E(n1041), .F(
        n1042), .Y(n1037) );
  OAI21X1 U445 ( .B(n1038), .C(n1043), .A(n1044), .Y(n1040) );
  NOR3XL U446 ( .A(n1046), .B(n1042), .C(n2016), .Y(n1039) );
  NAND4X1 U447 ( .A(n2016), .B(n1038), .C(n1043), .D(n1045), .Y(n1044) );
  INVX1 U448 ( .A(n891), .Y(n2085) );
  NAND21X1 U449 ( .B(n446), .A(n15), .Y(n2087) );
  AOI21BBXL U450 ( .B(n1896), .C(n1730), .A(n1708), .Y(n1706) );
  NAND32X1 U451 ( .B(n529), .C(n521), .A(n1227), .Y(n524) );
  NAND21X1 U452 ( .B(n1898), .A(n877), .Y(n957) );
  INVX1 U453 ( .A(n999), .Y(n1911) );
  AO21X1 U454 ( .B(n1434), .C(n1415), .A(n1414), .Y(n1416) );
  GEN2XL U455 ( .D(n1413), .E(n660), .C(n1523), .B(n176), .A(n1412), .Y(n1414)
         );
  AOI31X1 U456 ( .A(n1411), .B(n1587), .C(n1410), .D(n1413), .Y(n1412) );
  NOR3XL U457 ( .A(n1730), .B(n90), .C(n1708), .Y(n1707) );
  NAND2X1 U458 ( .A(n1593), .B(n1911), .Y(n917) );
  INVX1 U459 ( .A(n892), .Y(n2092) );
  INVX1 U460 ( .A(n528), .Y(n1929) );
  INVX1 U461 ( .A(n444), .Y(n442) );
  INVX1 U462 ( .A(n375), .Y(n377) );
  INVX1 U463 ( .A(n375), .Y(n380) );
  INVX1 U464 ( .A(n375), .Y(n376) );
  NOR3XL U465 ( .A(n2092), .B(n2097), .C(n2030), .Y(n1731) );
  INVX1 U466 ( .A(n1167), .Y(n2042) );
  INVX1 U467 ( .A(n1185), .Y(n2046) );
  INVX1 U468 ( .A(n1773), .Y(n1841) );
  NAND21X1 U469 ( .B(n430), .A(n1670), .Y(n1456) );
  NAND21X1 U470 ( .B(n2100), .A(n1948), .Y(n2037) );
  NAND21X1 U471 ( .B(n1274), .A(n725), .Y(n1971) );
  OR2X1 U472 ( .A(n528), .B(n1508), .Y(n488) );
  NAND21X1 U473 ( .B(n429), .A(n946), .Y(n658) );
  INVX1 U474 ( .A(n2039), .Y(n1948) );
  NAND32X1 U475 ( .B(n1291), .C(n397), .A(n1885), .Y(n678) );
  INVX1 U476 ( .A(n2088), .Y(n1922) );
  INVX1 U477 ( .A(n2044), .Y(n1921) );
  INVX1 U478 ( .A(n1176), .Y(n1926) );
  INVX1 U479 ( .A(n815), .Y(n1896) );
  INVX1 U480 ( .A(n369), .Y(n372) );
  INVX1 U481 ( .A(n369), .Y(n371) );
  INVX1 U482 ( .A(n369), .Y(n373) );
  INVX1 U483 ( .A(n2043), .Y(n946) );
  INVX1 U484 ( .A(n604), .Y(n1917) );
  AND3X1 U485 ( .A(N11493), .B(codefetch_s), .C(n1886), .Y(N671) );
  NAND2X1 U486 ( .A(n1179), .B(n1186), .Y(n1200) );
  OAI32X1 U487 ( .A(codefetch_s), .B(n721), .C(n695), .D(n722), .E(n1274), .Y(
        N679) );
  INVX1 U488 ( .A(n445), .Y(n370) );
  INVX1 U489 ( .A(n964), .Y(n1913) );
  OR2X1 U490 ( .A(n722), .B(n1971), .Y(n727) );
  NAND2X1 U491 ( .A(n2080), .B(n1947), .Y(n1726) );
  NAND2X1 U492 ( .A(n1726), .B(n1680), .Y(n1156) );
  OAI31XL U493 ( .A(n1997), .B(n1971), .C(n399), .D(n720), .Y(N675) );
  OAI31XL U494 ( .A(n1971), .B(n1999), .C(n399), .D(n720), .Y(N677) );
  INVX1 U495 ( .A(n1365), .Y(n2047) );
  INVX1 U496 ( .A(ramdatai[5]), .Y(n2169) );
  INVX1 U497 ( .A(ramdatai[4]), .Y(n2170) );
  INVX1 U498 ( .A(ramdatai[6]), .Y(n2168) );
  OAI21BBX1 U499 ( .A(n1886), .B(N11494), .C(n720), .Y(N672) );
  OAI21BBX1 U500 ( .A(n1886), .B(N11492), .C(n720), .Y(N670) );
  INVX1 U501 ( .A(n1043), .Y(n1990) );
  INVX1 U502 ( .A(n1119), .Y(n2082) );
  INVX1 U503 ( .A(ramdatai[7]), .Y(n2167) );
  INVX1 U504 ( .A(ramdatai[3]), .Y(n2171) );
  INVX1 U505 ( .A(ramdatai[2]), .Y(n2172) );
  NAND21X1 U506 ( .B(n429), .A(n168), .Y(n668) );
  AO21X1 U507 ( .B(n1227), .C(n529), .A(n769), .Y(n608) );
  AO21X1 U508 ( .B(n568), .C(n1016), .A(n2077), .Y(n628) );
  INVX1 U509 ( .A(n908), .Y(n568) );
  NAND32X1 U510 ( .B(n519), .C(n529), .A(n521), .Y(n1196) );
  OR2X1 U511 ( .A(n430), .B(n1582), .Y(n690) );
  AO21X1 U512 ( .B(n1118), .C(n1946), .A(n1605), .Y(n1344) );
  AND2X1 U513 ( .A(n1489), .B(n1911), .Y(n1609) );
  NAND5XL U514 ( .A(n169), .B(n1908), .C(n655), .D(n170), .E(n668), .Y(n651)
         );
  NAND21X1 U515 ( .B(n1583), .A(n2035), .Y(n572) );
  NAND21X1 U516 ( .B(n1159), .A(n576), .Y(n1580) );
  NAND32X1 U517 ( .B(n999), .C(n583), .A(n1907), .Y(n1577) );
  NAND21X1 U518 ( .B(n1159), .A(n992), .Y(n1578) );
  NAND21X1 U519 ( .B(n1159), .A(n1021), .Y(n1586) );
  INVX1 U520 ( .A(n1159), .Y(n1907) );
  INVX1 U521 ( .A(n560), .Y(n1919) );
  INVX1 U522 ( .A(n1032), .Y(n2070) );
  INVX1 U523 ( .A(n1227), .Y(n519) );
  NAND2X1 U524 ( .A(n2050), .B(n1647), .Y(n1363) );
  NAND2X1 U525 ( .A(n2049), .B(n1647), .Y(n1364) );
  NOR3XL U526 ( .A(n2100), .B(n2042), .C(n917), .Y(n1583) );
  AND2X1 U527 ( .A(n401), .B(n1075), .Y(N588) );
  NOR2X1 U528 ( .A(n2101), .B(n2097), .Y(n1737) );
  INVX1 U529 ( .A(n571), .Y(n576) );
  NAND21X1 U530 ( .B(instr[5]), .A(n1673), .Y(n571) );
  INVX1 U531 ( .A(n432), .Y(n430) );
  INVX1 U532 ( .A(n432), .Y(n431) );
  INVX1 U533 ( .A(n1116), .Y(n2095) );
  INVX1 U534 ( .A(n629), .Y(n624) );
  OR2X1 U535 ( .A(n430), .B(n1581), .Y(n666) );
  INVX1 U536 ( .A(n720), .Y(n1972) );
  NAND2X1 U537 ( .A(n1608), .B(n972), .Y(n978) );
  INVX1 U538 ( .A(N11528), .Y(n2109) );
  NAND2X1 U539 ( .A(n1737), .B(n892), .Y(n1600) );
  INVX1 U540 ( .A(n646), .Y(n655) );
  INVX1 U541 ( .A(n1599), .Y(n583) );
  INVX1 U542 ( .A(n1704), .Y(n713) );
  INVX1 U543 ( .A(n1705), .Y(n710) );
  INVX1 U544 ( .A(n1597), .Y(n575) );
  NAND21X1 U545 ( .B(n170), .A(n645), .Y(n1572) );
  NAND21X1 U546 ( .B(n601), .A(n772), .Y(n1158) );
  NAND21X1 U547 ( .B(n612), .A(n777), .Y(n614) );
  NAND21X1 U548 ( .B(n770), .A(n1666), .Y(n590) );
  OR2X1 U549 ( .A(n538), .B(n536), .Y(n1470) );
  INVX1 U550 ( .A(n1515), .Y(n1904) );
  NOR2X1 U551 ( .A(n2029), .B(n2083), .Y(n909) );
  NOR2X1 U552 ( .A(n9), .B(n446), .Y(n1061) );
  INVX1 U553 ( .A(n618), .Y(n619) );
  INVX1 U554 ( .A(n617), .Y(n621) );
  NAND21X1 U555 ( .B(n620), .A(n618), .Y(n617) );
  INVX1 U556 ( .A(n1422), .Y(n1537) );
  INVX1 U557 ( .A(n578), .Y(n645) );
  NAND21X1 U558 ( .B(n646), .A(n654), .Y(n578) );
  INVX1 U559 ( .A(n1494), .Y(n555) );
  INVX1 U560 ( .A(n541), .Y(n770) );
  NAND2X1 U561 ( .A(n1112), .B(n2085), .Y(n1857) );
  INVX1 U562 ( .A(n916), .Y(n2041) );
  NAND21X1 U563 ( .B(n169), .A(n645), .Y(n1584) );
  NAND31X1 U564 ( .C(n635), .A(n1611), .B(n930), .Y(n1458) );
  NAND21X1 U565 ( .B(n150), .A(n972), .Y(n921) );
  NAND21X1 U566 ( .B(n2099), .A(n891), .Y(n809) );
  OR2X1 U567 ( .A(instr[5]), .B(n612), .Y(n811) );
  NAND32X1 U568 ( .B(n921), .C(n792), .A(n791), .Y(n1759) );
  NOR43XL U569 ( .B(n1581), .C(n1847), .D(n1582), .A(n1583), .Y(n717) );
  NOR43XL U570 ( .B(n1580), .C(n1578), .D(n1586), .A(n168), .Y(n1847) );
  OAI21X1 U571 ( .B(n2029), .C(n2084), .A(n1638), .Y(n922) );
  NAND31X1 U572 ( .C(n909), .A(n2035), .B(n1680), .Y(n1677) );
  NOR2X1 U573 ( .A(n2101), .B(n2095), .Y(n1686) );
  XNOR2XL U574 ( .A(n983), .B(n1086), .Y(n556) );
  AO21X1 U575 ( .B(n1609), .C(n15), .A(n977), .Y(n627) );
  NOR2X1 U576 ( .A(n2096), .B(n9), .Y(n1640) );
  INVX1 U577 ( .A(n960), .Y(n950) );
  INVX1 U578 ( .A(n603), .Y(n808) );
  AND2X1 U579 ( .A(n1834), .B(n1922), .Y(n1798) );
  INVX1 U580 ( .A(n635), .Y(n644) );
  OR3XL U581 ( .A(n1799), .B(n1798), .C(n1793), .Y(n1833) );
  INVX1 U582 ( .A(n2035), .Y(n782) );
  INVX1 U583 ( .A(n2096), .Y(n1892) );
  INVX1 U584 ( .A(n632), .Y(n1910) );
  NOR2X1 U585 ( .A(n2088), .B(n916), .Y(n1799) );
  OAI21X1 U586 ( .B(n2097), .C(n2030), .A(n1871), .Y(n1873) );
  NOR2X1 U587 ( .A(n2029), .B(n2088), .Y(n1794) );
  INVX1 U588 ( .A(n1634), .Y(n386) );
  NOR4XL U589 ( .A(n918), .B(n919), .C(n920), .D(n921), .Y(n905) );
  NAND3X1 U590 ( .A(n1577), .B(n1579), .C(n1585), .Y(n924) );
  NOR2X1 U591 ( .A(n2029), .B(n2092), .Y(n1789) );
  NAND3X1 U592 ( .A(n1829), .B(n1830), .C(n1831), .Y(n920) );
  NOR43XL U593 ( .B(n1760), .C(n1166), .D(n1758), .A(n1772), .Y(n1830) );
  NOR4XL U594 ( .A(n1888), .B(n1887), .C(n1786), .D(n1787), .Y(n1829) );
  NOR4XL U595 ( .A(n1832), .B(n1833), .C(n1794), .D(n1782), .Y(n1831) );
  NAND4X1 U596 ( .A(n1771), .B(n1777), .C(n1776), .D(n1781), .Y(n1832) );
  NAND3X1 U597 ( .A(n2043), .B(n897), .C(n898), .Y(n750) );
  INVX1 U598 ( .A(n1759), .Y(n898) );
  INVX1 U599 ( .A(n1331), .Y(n2099) );
  OR3XL U600 ( .A(n1788), .B(n1640), .C(n1789), .Y(n150) );
  NAND21X1 U601 ( .B(n1159), .A(n1017), .Y(n1166) );
  NAND32X1 U602 ( .B(n1159), .C(n583), .A(n960), .Y(n716) );
  INVX1 U603 ( .A(n601), .Y(n1022) );
  INVX1 U604 ( .A(n656), .Y(n657) );
  NOR2X1 U605 ( .A(n916), .B(n2083), .Y(n1772) );
  INVX1 U606 ( .A(n581), .Y(n636) );
  NAND21X1 U607 ( .B(n1611), .A(n930), .Y(n581) );
  NOR2X1 U608 ( .A(n2030), .B(n2100), .Y(n915) );
  INVX1 U609 ( .A(n1533), .Y(n2014) );
  INVX1 U610 ( .A(n865), .Y(n2015) );
  INVX1 U611 ( .A(n853), .Y(n2013) );
  INVX1 U612 ( .A(n847), .Y(n2012) );
  INVX1 U613 ( .A(n841), .Y(n2011) );
  INVX1 U614 ( .A(n994), .Y(n1887) );
  NAND21X1 U615 ( .B(n960), .A(n1022), .Y(n994) );
  NAND3X1 U616 ( .A(n4), .B(n1639), .C(n1608), .Y(n918) );
  INVX1 U617 ( .A(n1683), .Y(n2084) );
  NAND2X1 U618 ( .A(n1686), .B(n892), .Y(n885) );
  NAND21X1 U619 ( .B(n999), .A(n1022), .Y(n949) );
  NAND21X1 U620 ( .B(n1159), .A(n1948), .Y(n796) );
  INVX1 U621 ( .A(n791), .Y(n910) );
  OAI21X1 U622 ( .B(n369), .C(n2102), .A(n2101), .Y(n894) );
  OAI22X1 U623 ( .A(n916), .B(n2084), .C(n2083), .D(n2094), .Y(n914) );
  NAND21X1 U624 ( .B(n382), .A(n1904), .Y(n1444) );
  INVX1 U625 ( .A(n2002), .Y(n1932) );
  INVX1 U626 ( .A(n2004), .Y(n1934) );
  INVX1 U627 ( .A(n2003), .Y(n1933) );
  INVX1 U628 ( .A(n2005), .Y(n1935) );
  INVX1 U629 ( .A(n2006), .Y(n1936) );
  INVX1 U630 ( .A(n2001), .Y(n1931) );
  INVX1 U631 ( .A(n2007), .Y(n1937) );
  NAND21X1 U632 ( .B(n1641), .A(n181), .Y(n1256) );
  NAND21X1 U633 ( .B(n1641), .A(n179), .Y(n1254) );
  NAND21X1 U634 ( .B(n1641), .A(n178), .Y(n1252) );
  NAND21X1 U635 ( .B(n1641), .A(n180), .Y(n1250) );
  NAND21X1 U636 ( .B(n1898), .A(n833), .Y(n818) );
  NAND21X1 U637 ( .B(n2017), .A(n389), .Y(n997) );
  INVX1 U638 ( .A(n490), .Y(n504) );
  NAND21X1 U639 ( .B(n491), .A(n1348), .Y(n490) );
  NAND21X1 U640 ( .B(n1610), .A(n387), .Y(n1342) );
  NAND21X1 U641 ( .B(n1949), .A(n388), .Y(n491) );
  NAND2X1 U642 ( .A(n1244), .B(n387), .Y(n1242) );
  NAND21X1 U643 ( .B(n1808), .A(n1168), .Y(n1170) );
  NAND21X1 U644 ( .B(n725), .A(n388), .Y(n721) );
  AO21X1 U645 ( .B(n395), .C(n484), .A(n462), .Y(N12697) );
  INVX1 U646 ( .A(n1241), .Y(n484) );
  AO21X1 U647 ( .B(n395), .C(n944), .A(n462), .Y(N12699) );
  INVX1 U648 ( .A(n1239), .Y(n944) );
  AO21X1 U649 ( .B(n395), .C(n945), .A(n462), .Y(N12698) );
  INVX1 U650 ( .A(n1240), .Y(n945) );
  AO21X1 U651 ( .B(n395), .C(n180), .A(n461), .Y(N12556) );
  AO21X1 U652 ( .B(n395), .C(n179), .A(n461), .Y(N12538) );
  AO21X1 U653 ( .B(n395), .C(n178), .A(n462), .Y(N12547) );
  AO21X1 U654 ( .B(n395), .C(n181), .A(n462), .Y(N12529) );
  INVX1 U655 ( .A(n837), .Y(n1898) );
  NOR2X1 U656 ( .A(n1158), .B(n429), .Y(n1307) );
  AND2X1 U657 ( .A(n1939), .B(n730), .Y(N583) );
  NAND2X1 U658 ( .A(n1007), .B(n1944), .Y(n1001) );
  OAI22X1 U659 ( .A(n1168), .B(n2000), .C(n158), .D(n1170), .Y(N12705) );
  OAI22X1 U660 ( .A(n817), .B(n93), .C(n1981), .D(n1264), .Y(N12494) );
  OAI22X1 U661 ( .A(n817), .B(n108), .C(n1981), .D(n1262), .Y(N12503) );
  OAI22X1 U662 ( .A(n817), .B(n81), .C(n1981), .D(n1260), .Y(N12512) );
  OAI22X1 U663 ( .A(n817), .B(n72), .C(n1981), .D(n1258), .Y(N12521) );
  OAI22X1 U664 ( .A(n817), .B(n84), .C(n1981), .D(n1256), .Y(N12530) );
  OAI22X1 U665 ( .A(n817), .B(n95), .C(n1981), .D(n1254), .Y(N12539) );
  OAI22X1 U666 ( .A(n817), .B(n67), .C(n1981), .D(n1252), .Y(N12548) );
  OAI22X1 U667 ( .A(n817), .B(n74), .C(n1981), .D(n1250), .Y(N12557) );
  OAI22X1 U668 ( .A(n872), .B(n84), .C(n1988), .D(n1256), .Y(N12603) );
  OAI22X1 U669 ( .A(n866), .B(n84), .C(n1987), .D(n1256), .Y(N12604) );
  OAI22X1 U670 ( .A(n860), .B(n84), .C(n1986), .D(n1256), .Y(N12605) );
  OAI22X1 U671 ( .A(n854), .B(n84), .C(n1985), .D(n1256), .Y(N12606) );
  OAI22X1 U672 ( .A(n842), .B(n84), .C(n1983), .D(n1256), .Y(N12608) );
  OAI22X1 U673 ( .A(n836), .B(n84), .C(n1982), .D(n1256), .Y(N12609) );
  OAI22X1 U674 ( .A(n812), .B(n84), .C(n1980), .D(n1256), .Y(N12531) );
  OAI22X1 U675 ( .A(n872), .B(n95), .C(n1988), .D(n1254), .Y(N12612) );
  OAI22X1 U676 ( .A(n866), .B(n95), .C(n1987), .D(n1254), .Y(N12613) );
  OAI22X1 U677 ( .A(n860), .B(n95), .C(n1986), .D(n1254), .Y(N12614) );
  OAI22X1 U678 ( .A(n854), .B(n95), .C(n1985), .D(n1254), .Y(N12615) );
  OAI22X1 U679 ( .A(n842), .B(n95), .C(n1983), .D(n1254), .Y(N12617) );
  OAI22X1 U680 ( .A(n836), .B(n95), .C(n1982), .D(n1254), .Y(N12618) );
  OAI22X1 U681 ( .A(n812), .B(n95), .C(n1980), .D(n1254), .Y(N12540) );
  OAI22X1 U682 ( .A(n872), .B(n67), .C(n1988), .D(n1252), .Y(N12621) );
  OAI22X1 U683 ( .A(n866), .B(n67), .C(n1987), .D(n1252), .Y(N12622) );
  OAI22X1 U684 ( .A(n860), .B(n67), .C(n1986), .D(n1252), .Y(N12623) );
  OAI22X1 U685 ( .A(n854), .B(n67), .C(n1985), .D(n1252), .Y(N12624) );
  OAI22X1 U686 ( .A(n842), .B(n67), .C(n1983), .D(n1252), .Y(N12626) );
  OAI22X1 U687 ( .A(n836), .B(n67), .C(n1982), .D(n1252), .Y(N12627) );
  OAI22X1 U688 ( .A(n812), .B(n67), .C(n1980), .D(n1252), .Y(N12549) );
  OAI22X1 U689 ( .A(n872), .B(n74), .C(n1988), .D(n1250), .Y(N12630) );
  OAI22X1 U690 ( .A(n866), .B(n74), .C(n1987), .D(n1250), .Y(N12631) );
  OAI22X1 U691 ( .A(n860), .B(n74), .C(n1986), .D(n1250), .Y(N12632) );
  OAI22X1 U692 ( .A(n854), .B(n74), .C(n1985), .D(n1250), .Y(N12633) );
  OAI22X1 U693 ( .A(n842), .B(n74), .C(n1983), .D(n1250), .Y(N12635) );
  OAI22X1 U694 ( .A(n836), .B(n74), .C(n1982), .D(n1250), .Y(N12636) );
  OAI22X1 U695 ( .A(n812), .B(n74), .C(n1980), .D(n1250), .Y(N12558) );
  OAI22X1 U696 ( .A(n872), .B(n93), .C(n1988), .D(n1264), .Y(N12567) );
  OAI22X1 U697 ( .A(n866), .B(n93), .C(n1987), .D(n1264), .Y(N12568) );
  OAI22X1 U698 ( .A(n860), .B(n93), .C(n1986), .D(n1264), .Y(N12569) );
  OAI22X1 U699 ( .A(n854), .B(n93), .C(n1985), .D(n1264), .Y(N12570) );
  OAI22X1 U700 ( .A(n842), .B(n93), .C(n1983), .D(n1264), .Y(N12572) );
  OAI22X1 U701 ( .A(n836), .B(n93), .C(n1982), .D(n1264), .Y(N12573) );
  OAI22X1 U702 ( .A(n812), .B(n93), .C(n1980), .D(n1264), .Y(N12495) );
  OAI22X1 U703 ( .A(n872), .B(n108), .C(n1988), .D(n1262), .Y(N12576) );
  OAI22X1 U704 ( .A(n866), .B(n108), .C(n1987), .D(n1262), .Y(N12577) );
  OAI22X1 U705 ( .A(n860), .B(n108), .C(n1986), .D(n1262), .Y(N12578) );
  OAI22X1 U706 ( .A(n854), .B(n108), .C(n1985), .D(n1262), .Y(N12579) );
  OAI22X1 U707 ( .A(n842), .B(n108), .C(n1983), .D(n1262), .Y(N12581) );
  OAI22X1 U708 ( .A(n836), .B(n108), .C(n1982), .D(n1262), .Y(N12582) );
  OAI22X1 U709 ( .A(n812), .B(n108), .C(n1980), .D(n1262), .Y(N12504) );
  OAI22X1 U710 ( .A(n872), .B(n81), .C(n1988), .D(n1260), .Y(N12585) );
  OAI22X1 U711 ( .A(n866), .B(n81), .C(n1987), .D(n1260), .Y(N12586) );
  OAI22X1 U712 ( .A(n860), .B(n81), .C(n1986), .D(n1260), .Y(N12587) );
  OAI22X1 U713 ( .A(n854), .B(n81), .C(n1985), .D(n1260), .Y(N12588) );
  OAI22X1 U714 ( .A(n842), .B(n81), .C(n1983), .D(n1260), .Y(N12590) );
  OAI22X1 U715 ( .A(n836), .B(n81), .C(n1982), .D(n1260), .Y(N12591) );
  OAI22X1 U716 ( .A(n812), .B(n81), .C(n1980), .D(n1260), .Y(N12513) );
  OAI22X1 U717 ( .A(n872), .B(n72), .C(n1988), .D(n1258), .Y(N12594) );
  OAI22X1 U718 ( .A(n866), .B(n72), .C(n1987), .D(n1258), .Y(N12595) );
  OAI22X1 U719 ( .A(n860), .B(n72), .C(n1986), .D(n1258), .Y(N12596) );
  OAI22X1 U720 ( .A(n854), .B(n72), .C(n1985), .D(n1258), .Y(N12597) );
  OAI22X1 U721 ( .A(n842), .B(n72), .C(n1983), .D(n1258), .Y(N12599) );
  OAI22X1 U722 ( .A(n836), .B(n72), .C(n1982), .D(n1258), .Y(N12600) );
  OAI22X1 U723 ( .A(n812), .B(n72), .C(n1980), .D(n1258), .Y(N12522) );
  OAI21X1 U724 ( .B(n1000), .C(n1001), .A(n453), .Y(N13293) );
  OAI21X1 U725 ( .B(n2073), .C(n1001), .A(n453), .Y(N13275) );
  OAI21X1 U726 ( .B(n1661), .C(n1001), .A(n453), .Y(N13266) );
  OAI21X1 U727 ( .B(n1000), .C(n1009), .A(n453), .Y(N13221) );
  OAI21X1 U728 ( .B(n2073), .C(n1009), .A(n453), .Y(N13203) );
  OAI21X1 U729 ( .B(n1661), .C(n1009), .A(n454), .Y(N13194) );
  OAI21X1 U730 ( .B(n1000), .C(n1011), .A(n454), .Y(N13149) );
  OAI21X1 U731 ( .B(n2073), .C(n1011), .A(n454), .Y(N13131) );
  OAI21X1 U732 ( .B(n1661), .C(n1011), .A(n454), .Y(N13122) );
  OAI31XL U733 ( .A(n1245), .B(dps[1]), .C(dps[0]), .D(n457), .Y(N12665) );
  OAI31XL U734 ( .A(n1247), .B(dps[1]), .C(dps[0]), .D(n463), .Y(N12637) );
  INVX1 U735 ( .A(n2000), .Y(n1930) );
  NAND2X1 U736 ( .A(n1246), .B(dps[2]), .Y(n1245) );
  NAND2X1 U737 ( .A(n452), .B(n2002), .Y(N12692) );
  NAND2X1 U738 ( .A(n452), .B(n2004), .Y(N12690) );
  NAND2X1 U739 ( .A(n452), .B(n2003), .Y(N12691) );
  OAI211X1 U740 ( .C(n695), .D(n721), .A(n722), .B(n456), .Y(N685) );
  INVX1 U741 ( .A(n1028), .Y(N10579) );
  NAND21X1 U742 ( .B(n1765), .A(n389), .Y(n1028) );
  INVX1 U743 ( .A(n1665), .Y(n1243) );
  NAND21X1 U744 ( .B(n1244), .A(n387), .Y(n1665) );
  AND2X1 U745 ( .A(n394), .B(n151), .Y(N10575) );
  NAND4X1 U746 ( .A(n1774), .B(n1775), .C(n1776), .D(n1777), .Y(n151) );
  NOR21XL U747 ( .B(n394), .A(n1783), .Y(N10573) );
  NOR4XL U748 ( .A(n1784), .B(n1785), .C(n1786), .D(n1787), .Y(n1783) );
  NOR21XL U749 ( .B(n394), .A(n1790), .Y(N10571) );
  NOR4XL U750 ( .A(n1791), .B(n1792), .C(n1793), .D(n1794), .Y(n1790) );
  NOR21XL U751 ( .B(n394), .A(n1768), .Y(N10576) );
  NOR43XL U752 ( .B(n1769), .C(n1770), .D(n1771), .A(n1772), .Y(n1768) );
  NOR21XL U753 ( .B(n394), .A(n1795), .Y(N10570) );
  NOR4XL U754 ( .A(n1796), .B(n1797), .C(n1798), .D(n1799), .Y(n1795) );
  NOR21XL U755 ( .B(n394), .A(n1778), .Y(N10574) );
  NOR43XL U756 ( .B(n1779), .C(n1780), .D(n1781), .A(n1782), .Y(n1778) );
  NAND21X1 U757 ( .B(n1808), .A(n1515), .Y(n1382) );
  INVX1 U758 ( .A(n486), .Y(n500) );
  AND2X1 U759 ( .A(n392), .B(n114), .Y(N12709) );
  AND2X1 U760 ( .A(n391), .B(n1455), .Y(N11485) );
  AND2X1 U761 ( .A(n500), .B(n493), .Y(N13372) );
  AND2X1 U762 ( .A(n500), .B(n494), .Y(N13370) );
  AND2X1 U763 ( .A(n500), .B(n495), .Y(N13368) );
  AND2X1 U764 ( .A(n500), .B(n496), .Y(N13373) );
  AND2X1 U765 ( .A(n500), .B(n497), .Y(N13371) );
  AND2X1 U766 ( .A(n500), .B(n498), .Y(N13369) );
  AND2X1 U767 ( .A(n1889), .B(n393), .Y(N10581) );
  AND2X1 U768 ( .A(n1888), .B(n392), .Y(N10586) );
  AND2X1 U769 ( .A(n392), .B(n2066), .Y(N12710) );
  NOR21XL U770 ( .B(n392), .A(n1236), .Y(N12702) );
  NOR21XL U771 ( .B(n391), .A(n1237), .Y(N12701) );
  NOR21XL U772 ( .B(n392), .A(n1235), .Y(N12703) );
  NOR21XL U773 ( .B(n391), .A(n1238), .Y(N12700) );
  AND2X1 U774 ( .A(n391), .B(n166), .Y(N12704) );
  AND2X1 U775 ( .A(n391), .B(sfrwe_comb_s), .Y(N11489) );
  AND2X1 U776 ( .A(n390), .B(n156), .Y(N11480) );
  AND2X1 U777 ( .A(n1766), .B(n392), .Y(N10578) );
  AND2X1 U778 ( .A(n390), .B(n157), .Y(N11479) );
  NOR21XL U779 ( .B(n390), .A(n1803), .Y(N10566) );
  NOR21XL U780 ( .B(n390), .A(n1760), .Y(N10584) );
  NOR21XL U781 ( .B(n401), .A(n1758), .Y(N10587) );
  AND2X1 U782 ( .A(n401), .B(n1451), .Y(N11478) );
  NOR2X1 U783 ( .A(n429), .B(n723), .Y(N681) );
  INVX1 U784 ( .A(n696), .Y(n1248) );
  INVX1 U785 ( .A(n970), .Y(n828) );
  INVX1 U786 ( .A(n1539), .Y(n1362) );
  MUX2X1 U787 ( .D0(n1576), .D1(n1584), .S(n1603), .Y(n1588) );
  MUX2X1 U788 ( .D0(n1584), .D1(n1576), .S(n176), .Y(n1410) );
  INVX1 U789 ( .A(n1511), .Y(n1914) );
  INVX1 U790 ( .A(n1512), .Y(n1924) );
  INVX1 U791 ( .A(n1510), .Y(n1915) );
  NAND2X1 U792 ( .A(n1467), .B(n1468), .Y(n1391) );
  INVX1 U793 ( .A(n5), .Y(n1587) );
  MUX2X1 U794 ( .D0(n1584), .D1(n1576), .S(n177), .Y(n1420) );
  INVX1 U795 ( .A(n1457), .Y(n1906) );
  ENOX1 U796 ( .A(n871), .B(n2090), .C(n964), .D(n1070), .Y(n1098) );
  INVX1 U797 ( .A(n1424), .Y(n1950) );
  NAND2X1 U798 ( .A(n2080), .B(n1489), .Y(n1468) );
  AND2X1 U799 ( .A(n1938), .B(n2072), .Y(n742) );
  NOR2X1 U800 ( .A(n1325), .B(n1244), .Y(n1271) );
  NOR2X1 U801 ( .A(n1327), .B(n1244), .Y(n1269) );
  NOR2X1 U802 ( .A(n1326), .B(n1244), .Y(n1270) );
  NAND2X1 U803 ( .A(n2040), .B(n1129), .Y(n1153) );
  NOR21XL U804 ( .B(n1328), .A(n1244), .Y(n1267) );
  NAND4X1 U805 ( .A(n1327), .B(n1329), .C(n1325), .D(n1326), .Y(n1328) );
  INVX1 U806 ( .A(n1089), .Y(n2027) );
  NAND2X1 U807 ( .A(n1105), .B(n1106), .Y(n1068) );
  NOR2X1 U808 ( .A(n1125), .B(n429), .Y(n1072) );
  NAND41X1 U809 ( .D(n920), .A(n1806), .B(n1805), .C(n1827), .Y(n1826) );
  NOR32XL U810 ( .B(n1803), .C(n1802), .A(n1890), .Y(n1827) );
  NOR4XL U811 ( .A(n1823), .B(n1824), .C(n1825), .D(n1826), .Y(n1818) );
  NAND4X1 U812 ( .A(n1780), .B(n1779), .C(n1774), .D(n1838), .Y(n1823) );
  NAND4X1 U813 ( .A(n1769), .B(n1775), .C(n1770), .D(n1837), .Y(n1824) );
  NAND4X1 U814 ( .A(n1800), .B(n1767), .C(n1801), .D(n1836), .Y(n1825) );
  INVX1 U815 ( .A(n1134), .Y(n2023) );
  INVX1 U816 ( .A(n1138), .Y(n962) );
  OAI21X1 U817 ( .B(n431), .C(n2091), .A(n1107), .Y(n1106) );
  NOR2X1 U818 ( .A(n885), .B(n429), .Y(n1071) );
  NOR42XL U819 ( .C(n1761), .D(n1762), .A(n1889), .B(n1766), .Y(n1836) );
  NAND2X1 U820 ( .A(n1828), .B(n1952), .Y(n1761) );
  NAND2X1 U821 ( .A(n1828), .B(n2080), .Y(n1762) );
  NAND2X1 U822 ( .A(n1062), .B(n1922), .Y(n1802) );
  NAND2X1 U823 ( .A(n1062), .B(n892), .Y(n1756) );
  NAND2X1 U824 ( .A(n1108), .B(n2025), .Y(n1094) );
  AND3X1 U825 ( .A(n117), .B(n437), .C(n435), .Y(n152) );
  AND3X1 U826 ( .A(n435), .B(n117), .C(n436), .Y(n153) );
  AND3X1 U827 ( .A(n117), .B(n437), .C(n434), .Y(n154) );
  AND3X1 U828 ( .A(n434), .B(n117), .C(n436), .Y(n155) );
  INVX1 U829 ( .A(n1066), .Y(n2090) );
  NAND31X1 U830 ( .C(n999), .A(n1828), .B(n15), .Y(n1806) );
  INVX1 U831 ( .A(n1070), .Y(n1087) );
  AND2X1 U832 ( .A(n1118), .B(n1061), .Y(n1785) );
  NAND2X1 U833 ( .A(n1834), .B(n1946), .Y(n1801) );
  NAND2X1 U834 ( .A(n1834), .B(n1683), .Y(n1767) );
  NAND2X1 U835 ( .A(n1062), .B(n1946), .Y(n1805) );
  INVX1 U836 ( .A(n990), .Y(n1890) );
  NAND32X1 U837 ( .B(n917), .C(n56), .A(n912), .Y(n990) );
  NOR4XL U838 ( .A(n1796), .B(n1797), .C(n1791), .D(n1792), .Y(n1838) );
  NOR2X1 U839 ( .A(n2094), .B(n2088), .Y(n1791) );
  OR2X1 U840 ( .A(n897), .B(n2190), .Y(n1764) );
  NAND2X1 U841 ( .A(n1032), .B(n452), .Y(n1029) );
  INVX1 U842 ( .A(rst), .Y(n463) );
  MUX2BXL U843 ( .D0(mempswr), .D1(n1469), .S(n451), .Y(mempswr_comb) );
  NAND21X1 U844 ( .B(n2072), .A(n730), .Y(n1459) );
  XOR3X1 U845 ( .A(n1552), .B(n6), .C(n1353), .Y(n758) );
  INVX1 U846 ( .A(n1553), .Y(n702) );
  NAND21X1 U847 ( .B(n656), .A(n650), .Y(n700) );
  NAND32X1 U848 ( .B(n1065), .C(n1804), .A(n806), .Y(n959) );
  OAI211X1 U849 ( .C(n555), .D(n648), .A(n554), .B(n553), .Y(n1086) );
  OA22X1 U850 ( .A(n1131), .B(n1512), .C(n1467), .D(n1091), .Y(n554) );
  OA222X1 U851 ( .A(n1225), .B(n1511), .C(n965), .D(n1510), .E(n1991), .F(n552), .Y(n553) );
  NAND21X1 U852 ( .B(memack), .A(n468), .Y(n465) );
  INVX1 U853 ( .A(sfrdatai[0]), .Y(n965) );
  INVX2 U854 ( .A(n1304), .Y(n1530) );
  OAI32X1 U855 ( .A(n871), .B(n2127), .C(n1521), .D(n752), .E(n746), .Y(n753)
         );
  INVX1 U856 ( .A(n471), .Y(n469) );
  OA22X1 U857 ( .A(n2173), .B(n555), .C(n1467), .D(n1913), .Y(n540) );
  OA222X1 U858 ( .A(n871), .B(n1512), .C(n552), .D(n1992), .E(n1511), .F(n2126), .Y(n539) );
  MUX2X1 U859 ( .D0(ramsfraddr[2]), .D1(n156), .S(n451), .Y(ramsfraddr_comb[2]) );
  NAND31X1 U860 ( .C(n1721), .A(n1716), .B(n1715), .Y(n1701) );
  OAI222XL U861 ( .A(n1997), .B(n1712), .C(n1989), .D(n1701), .E(n1716), .F(
        n1993), .Y(n156) );
  NOR8XL U862 ( .A(n964), .B(n963), .C(n868), .D(n1361), .E(n970), .F(n969), 
        .G(n968), .H(n967), .Y(n779) );
  OAI22X1 U863 ( .A(n1700), .B(n1999), .C(n1701), .D(n1035), .Y(n1455) );
  OA222X1 U864 ( .A(N13353), .B(n1183), .C(n1966), .D(n1666), .E(n1227), .F(
        n2053), .Y(n548) );
  NAND21X1 U865 ( .B(n840), .A(n823), .Y(n1193) );
  AND2X1 U866 ( .A(n1715), .B(n1716), .Y(n1700) );
  OAI222XL U867 ( .A(n1716), .B(n1991), .C(n1701), .D(n2016), .E(n1712), .F(
        n1995), .Y(n1451) );
  OAI222XL U868 ( .A(n1996), .B(n1712), .C(n1990), .D(n1701), .E(n1716), .F(
        n1992), .Y(n157) );
  INVX1 U869 ( .A(n822), .Y(n823) );
  NAND21X1 U870 ( .B(n834), .A(n821), .Y(n822) );
  NOR2X1 U871 ( .A(n1662), .B(memdatai[7]), .Y(n1721) );
  NAND2X1 U872 ( .A(n1721), .B(n1716), .Y(n1712) );
  INVX1 U873 ( .A(n718), .Y(sfrwe_comb_s) );
  NAND21X1 U874 ( .B(n1298), .A(n1297), .Y(n718) );
  OR2X1 U875 ( .A(n1662), .B(n1999), .Y(n1715) );
  NAND2X1 U876 ( .A(n806), .B(n808), .Y(n1160) );
  NAND2X1 U877 ( .A(n834), .B(n821), .Y(n1202) );
  MUX2X1 U878 ( .D0(ramsfraddr[1]), .D1(n157), .S(n451), .Y(ramsfraddr_comb[1]) );
  MUX2X1 U879 ( .D0(ramsfraddr[0]), .D1(n1451), .S(n450), .Y(
        ramsfraddr_comb[0]) );
  NAND21X1 U880 ( .B(n1234), .A(n1233), .Y(n1476) );
  AO2222XL U881 ( .A(alu_out[0]), .B(n113), .C(n384), .D(n1642), .E(n1896), 
        .F(ramdatai[0]), .G(n1897), .H(n1149), .Y(n1234) );
  OA2222XL U882 ( .A(n1225), .B(n1202), .C(n1991), .D(n1198), .E(n1197), .F(
        n1193), .G(n37), .H(n1161), .Y(n1233) );
  INVX1 U883 ( .A(n1131), .Y(n1149) );
  NAND21X1 U884 ( .B(n989), .A(n988), .Y(n1477) );
  AO2222XL U885 ( .A(alu_out[1]), .B(n1160), .C(n384), .D(n1643), .E(n1897), 
        .F(n986), .G(n1896), .H(ramdatai[1]), .Y(n989) );
  OA2222XL U886 ( .A(n2126), .B(n1202), .C(n1992), .D(n1198), .E(n987), .F(
        n1193), .G(n43), .H(n1161), .Y(n988) );
  INVX1 U887 ( .A(n871), .Y(n986) );
  NAND21X1 U888 ( .B(n980), .A(n979), .Y(n1491) );
  OA2222XL U889 ( .A(n31), .B(n976), .C(n2129), .D(n975), .E(n2053), .F(n974), 
        .G(n2150), .H(n973), .Y(n979) );
  AO2222XL U890 ( .A(n1612), .B(n384), .C(n971), .D(pc_i[8]), .E(n1898), .F(
        instr[5]), .G(alu_out[8]), .H(n113), .Y(n980) );
  INVX1 U891 ( .A(n963), .Y(n1091) );
  OA222X1 U892 ( .A(n2173), .B(n192), .C(n871), .D(n1565), .E(n1352), .F(n1563), .Y(n1354) );
  OAI21BBX1 U893 ( .A(codefetch_s), .B(n1960), .C(n726), .Y(n1052) );
  AOI22X1 U894 ( .A(incdec_out[7]), .B(n1422), .C(pc_i[7]), .D(n1906), .Y(
        n1394) );
  NAND21X1 U895 ( .B(n1064), .A(n1060), .Y(n1075) );
  MUX2X1 U896 ( .D0(n763), .D1(n1840), .S(codefetch_s), .Y(n1064) );
  MUX2X1 U897 ( .D0(n1059), .D1(n1058), .S(n680), .Y(n1060) );
  OAI21BBX1 U898 ( .A(n2008), .B(n680), .C(n684), .Y(n763) );
  OAI22AX1 U899 ( .D(N11547), .C(n2177), .A(n2178), .B(n2109), .Y(N11560) );
  NOR21XL U900 ( .B(n2178), .A(N11528), .Y(n2177) );
  OAI222XL U901 ( .A(n670), .B(n1450), .C(n1443), .D(n1444), .E(n2136), .F(
        n451), .Y(ramdatao_comb[6]) );
  INVX1 U902 ( .A(n1057), .Y(n1443) );
  OAI222XL U903 ( .A(n667), .B(n1450), .C(n1970), .D(n1444), .E(n2130), .F(
        n2184), .Y(ramdatao_comb[7]) );
  NAND2X1 U904 ( .A(n1371), .B(n2115), .Y(n1381) );
  AOI22AXL U905 ( .A(n2180), .B(N11527), .D(n2181), .C(N11546), .Y(n2178) );
  NOR2X1 U906 ( .A(N11527), .B(n2180), .Y(n2181) );
  AOI22X1 U907 ( .A(incdec_out[6]), .B(n1422), .C(pc_i[6]), .D(n1906), .Y(
        n1429) );
  XOR3X1 U908 ( .A(n1552), .B(n165), .C(n1551), .Y(incdec_out[6]) );
  INVX1 U909 ( .A(n1567), .Y(n1551) );
  AND3X1 U910 ( .A(n159), .B(n160), .C(n771), .Y(n158) );
  OA22X1 U911 ( .A(n1203), .B(n2133), .C(n1204), .D(n1185), .Y(n159) );
  MUX2IX1 U912 ( .D0(n1201), .D1(n1217), .S(N11584), .Y(n160) );
  NAND43X1 U913 ( .B(n597), .C(n596), .D(n595), .A(n594), .Y(n970) );
  OAI22X1 U914 ( .A(n2133), .B(n1196), .C(n1356), .D(n1556), .Y(n595) );
  OAI22X1 U915 ( .A(n1183), .B(n2159), .C(n2130), .D(n1227), .Y(n596) );
  AO21X1 U916 ( .B(multemp2[1]), .C(n1926), .A(n1400), .Y(n597) );
  XNOR2XL U917 ( .A(n1369), .B(n1370), .Y(N11549) );
  NOR2X1 U918 ( .A(n1371), .B(n2133), .Y(n1369) );
  OAI222XL U919 ( .A(n671), .B(n1450), .C(n1442), .D(n1444), .E(n2141), .F(
        waitstaten), .Y(ramdatao_comb[5]) );
  INVX1 U920 ( .A(n1055), .Y(n1442) );
  AOI222XL U921 ( .A(incdec_out[5]), .B(n1422), .C(ramdatai[5]), .D(n2079), 
        .E(n968), .F(n1398), .Y(n1448) );
  XOR3X1 U922 ( .A(n1552), .B(n164), .C(n1546), .Y(incdec_out[5]) );
  INVX1 U923 ( .A(n1548), .Y(n1546) );
  OAI21X1 U924 ( .B(n1372), .C(n2126), .A(n2107), .Y(N11523) );
  NAND2X1 U925 ( .A(n1967), .B(n2127), .Y(n1378) );
  INVX1 U926 ( .A(n1379), .Y(n2110) );
  OA222X1 U927 ( .A(n1343), .B(n1563), .C(n865), .D(n1565), .E(n2172), .F(n192), .Y(n161) );
  NAND21X1 U928 ( .B(n840), .A(n845), .Y(n877) );
  OA222X1 U929 ( .A(n1903), .B(n1539), .C(n1538), .D(n1553), .E(n1537), .F(
        n1536), .Y(n1496) );
  XOR3X1 U930 ( .A(n1552), .B(n162), .C(n1542), .Y(n1536) );
  GEN2XL U931 ( .D(n1524), .E(n660), .C(n1523), .B(n175), .A(n1522), .Y(n1528)
         );
  OAI222XL U932 ( .A(n672), .B(n1450), .C(n1418), .D(n1444), .E(n2134), .F(
        n451), .Y(ramdatao_comb[4]) );
  INVX1 U933 ( .A(n1056), .Y(n1418) );
  AOI222XL U934 ( .A(incdec_out[4]), .B(n1422), .C(ramdatai[4]), .D(n2079), 
        .E(n967), .F(n1398), .Y(n1472) );
  XOR3X1 U935 ( .A(n1552), .B(n163), .C(n1543), .Y(incdec_out[4]) );
  INVX1 U936 ( .A(n1545), .Y(n1543) );
  XNOR2XL U937 ( .A(n2178), .B(n2179), .Y(adder_out[6]) );
  XNOR2XL U938 ( .A(N11547), .B(n2109), .Y(n2179) );
  NAND3X1 U939 ( .A(n1923), .B(n1963), .C(n1012), .Y(n1168) );
  NOR2X1 U940 ( .A(n2128), .B(n1340), .Y(n1338) );
  NAND3X1 U941 ( .A(n1012), .B(n1943), .C(n1014), .Y(n1340) );
  NAND3X1 U942 ( .A(n2119), .B(n2121), .C(n2071), .Y(n1000) );
  OAI22X1 U943 ( .A(n1339), .B(n438), .C(n1340), .D(n2053), .Y(N346) );
  AND2X1 U944 ( .A(n1336), .B(n1335), .Y(n1339) );
  INVX1 U945 ( .A(n508), .Y(n1923) );
  NAND32X1 U946 ( .B(n1000), .C(n1962), .A(n831), .Y(n508) );
  INVX1 U947 ( .A(n1663), .Y(n1943) );
  INVX1 U948 ( .A(N347), .Y(n435) );
  OA222X1 U949 ( .A(n1534), .B(n1563), .C(n1533), .D(n1565), .E(n2171), .F(
        n192), .Y(n162) );
  MUX2AXL U950 ( .D0(rn[4]), .D1(n2134), .S(n580), .Y(n853) );
  MUX2X1 U951 ( .D0(n338), .D1(n333), .S(n2066), .Y(rn[4]) );
  MUX4X1 U952 ( .D0(n337), .D1(n335), .D2(n336), .D3(n334), .S0(n2065), .S1(
        n101), .Y(n338) );
  MUX4X1 U953 ( .D0(n332), .D1(n330), .D2(n331), .D3(n329), .S0(n2065), .S1(
        n101), .Y(n333) );
  NAND32X1 U954 ( .B(n534), .C(n533), .A(n532), .Y(n964) );
  OAI22X1 U955 ( .A(n1227), .B(n2064), .C(n1356), .D(n783), .Y(n534) );
  OA222X1 U956 ( .A(n560), .B(n2159), .C(n1967), .D(n2048), .E(n545), .F(n531), 
        .Y(n532) );
  OAI211X1 U957 ( .C(n1549), .D(n2126), .A(n526), .B(n525), .Y(n533) );
  MUX2AXL U958 ( .D0(rn[3]), .D1(n2128), .S(n580), .Y(n1533) );
  MUX2X1 U959 ( .D0(n328), .D1(n323), .S(n2066), .Y(rn[3]) );
  MUX4X1 U960 ( .D0(n327), .D1(n325), .D2(n326), .D3(n324), .S0(n2065), .S1(
        n100), .Y(n328) );
  MUX4X1 U961 ( .D0(n322), .D1(n320), .D2(n321), .D3(n319), .S0(n2065), .S1(
        n100), .Y(n323) );
  OAI221X1 U962 ( .A(n1702), .B(n1533), .C(n1713), .D(n1189), .E(n1717), .Y(
        n1041) );
  OA222X1 U963 ( .A(n1238), .B(n1703), .C(n2132), .D(n1705), .E(n2152), .F(
        n1704), .Y(n1717) );
  NAND21X1 U964 ( .B(mempsack), .A(n470), .Y(n466) );
  OAI222XL U965 ( .A(n673), .B(n1450), .C(n1994), .D(n1444), .E(n2120), .F(
        n450), .Y(ramdatao_comb[2]) );
  OA22X1 U966 ( .A(N13343), .B(n1183), .C(n2154), .D(n1176), .Y(n525) );
  NAND21X1 U967 ( .B(n1736), .A(n903), .Y(n1747) );
  NOR2X1 U968 ( .A(n1955), .B(n448), .Y(n891) );
  OAI221X1 U969 ( .A(n853), .B(n1702), .C(n1188), .D(n1713), .E(n1714), .Y(
        n1045) );
  OA222X1 U970 ( .A(n1237), .B(n1703), .C(n2163), .D(n1705), .E(n2155), .F(
        n1704), .Y(n1714) );
  NOR2X1 U971 ( .A(n2105), .B(n2085), .Y(n1683) );
  NAND2X1 U972 ( .A(irq), .B(n881), .Y(n725) );
  INVX1 U973 ( .A(n1763), .Y(n881) );
  OAI222XL U974 ( .A(n1606), .B(n1604), .C(n1603), .D(n1596), .E(n1595), .F(
        n1592), .Y(n1397) );
  AND3X1 U975 ( .A(n1588), .B(n1587), .C(n196), .Y(n1592) );
  OA21XL U976 ( .B(n1584), .C(n1574), .A(n1572), .Y(n1596) );
  INVXL U977 ( .A(n1574), .Y(n1595) );
  INVX1 U978 ( .A(n840), .Y(n846) );
  OAI221X1 U979 ( .A(n1562), .B(n1604), .C(n1561), .D(n1560), .E(n1559), .Y(
        n1431) );
  AOI211X1 U980 ( .C(n660), .D(n1555), .A(n197), .B(n5), .Y(n1560) );
  AO21X1 U981 ( .B(n1558), .C(n1572), .A(n1557), .Y(n1559) );
  MUX2X1 U982 ( .D0(n1556), .D1(n1965), .S(n1571), .Y(n1555) );
  AOI221XL U983 ( .A(pc_i[2]), .B(n1906), .C(n1368), .D(n1422), .E(n1367), .Y(
        n1388) );
  AO21X1 U984 ( .B(n1362), .C(n1361), .A(n1520), .Y(n1367) );
  XOR3X1 U985 ( .A(n1552), .B(n161), .C(n1359), .Y(n1368) );
  OAI22X1 U986 ( .A(n1499), .B(n33), .C(n1950), .D(n27), .Y(n1520) );
  AOI221XL U987 ( .A(n1438), .B(n177), .C(n1434), .D(n1433), .E(n1449), .Y(
        n1439) );
  OAI222XL U988 ( .A(n1456), .B(n2158), .C(n1457), .D(n2061), .E(n1458), .F(
        n2056), .Y(n1449) );
  AO21X1 U989 ( .B(n1432), .C(n660), .A(n1523), .Y(n1438) );
  ENOX1 U990 ( .A(n667), .B(n1382), .C(n1904), .D(N12476), .Y(N11505) );
  OA222X1 U991 ( .A(n1541), .B(n1563), .C(n853), .D(n1565), .E(n2170), .F(n192), .Y(n163) );
  OA222X1 U992 ( .A(n1544), .B(n1563), .C(n847), .D(n1565), .E(n2169), .F(n192), .Y(n164) );
  AND2X1 U993 ( .A(n1295), .B(n452), .Y(N512) );
  AOI211X1 U994 ( .C(n660), .D(n1330), .A(n1303), .B(n197), .Y(n1308) );
  MUX2AXL U995 ( .D0(n2053), .D1(n1300), .S(waitstaten), .Y(ramdatao_comb[0])
         );
  MUX2AXL U996 ( .D0(n2064), .D1(n1301), .S(waitstaten), .Y(ramdatao_comb[1])
         );
  NAND32X1 U997 ( .B(n1963), .C(n509), .A(n1923), .Y(n1227) );
  OA2222XL U998 ( .A(n1702), .B(n847), .C(n1236), .D(n1703), .E(n2157), .F(
        n1704), .G(n1963), .H(n1705), .Y(n1038) );
  NAND21X1 U999 ( .B(instr[5]), .A(n1956), .Y(n999) );
  NAND21X1 U1000 ( .B(n1002), .A(n1942), .Y(n1709) );
  NAND32X1 U1001 ( .B(n1729), .C(n2028), .A(n1499), .Y(n1708) );
  MUX2AXL U1002 ( .D0(rn[6]), .D1(n2136), .S(n580), .Y(n841) );
  MUX2X1 U1003 ( .D0(n358), .D1(n353), .S(n2066), .Y(rn[6]) );
  MUX4X1 U1004 ( .D0(n357), .D1(n355), .D2(n356), .D3(n354), .S0(n114), .S1(
        n101), .Y(n358) );
  MUX4X1 U1005 ( .D0(n352), .D1(n350), .D2(n351), .D3(n349), .S0(n114), .S1(
        n101), .Y(n353) );
  MUX2AXL U1006 ( .D0(rn[0]), .D1(n2053), .S(n580), .Y(n1131) );
  MUX2X1 U1007 ( .D0(n298), .D1(n293), .S(n2066), .Y(rn[0]) );
  MUX4X1 U1008 ( .D0(n297), .D1(n295), .D2(n296), .D3(n294), .S0(n114), .S1(
        n101), .Y(n298) );
  MUX4X1 U1009 ( .D0(n292), .D1(n290), .D2(n291), .D3(n289), .S0(n2065), .S1(
        n101), .Y(n293) );
  OA2222XL U1010 ( .A(n1702), .B(n841), .C(n1235), .D(n1703), .E(n1965), .F(
        n1704), .G(n1962), .H(n1705), .Y(n1042) );
  MUX2AXL U1011 ( .D0(rn[1]), .D1(n2064), .S(n580), .Y(n871) );
  MUX2X1 U1012 ( .D0(n308), .D1(n303), .S(n2066), .Y(rn[1]) );
  MUX4X1 U1013 ( .D0(n307), .D1(n305), .D2(n306), .D3(n304), .S0(n2065), .S1(
        n100), .Y(n308) );
  MUX4X1 U1014 ( .D0(n302), .D1(n300), .D2(n301), .D3(n299), .S0(n2065), .S1(
        n100), .Y(n303) );
  AND3X1 U1015 ( .A(n1223), .B(n1660), .C(n1920), .Y(n1647) );
  NAND3X1 U1016 ( .A(n1647), .B(n1649), .C(n1648), .Y(n528) );
  AO21X1 U1017 ( .B(n7), .C(n470), .A(n1690), .Y(n472) );
  MUX2AXL U1018 ( .D0(rn[5]), .D1(n2141), .S(n580), .Y(n847) );
  MUX2X1 U1019 ( .D0(n348), .D1(n343), .S(n2066), .Y(rn[5]) );
  MUX4X1 U1020 ( .D0(n347), .D1(n345), .D2(n346), .D3(n344), .S0(n114), .S1(
        n101), .Y(n348) );
  MUX4X1 U1021 ( .D0(n342), .D1(n340), .D2(n341), .D3(n339), .S0(n114), .S1(
        n101), .Y(n343) );
  OAI221X1 U1022 ( .A(n871), .B(n1702), .C(n1713), .D(n69), .E(n1720), .Y(
        n1043) );
  OA222X1 U1023 ( .A(n1240), .B(n1703), .C(n2119), .D(n1705), .E(n2151), .F(
        n1704), .Y(n1720) );
  INVX1 U1024 ( .A(n478), .Y(n1942) );
  NAND21X1 U1025 ( .B(n1663), .A(n1944), .Y(n478) );
  AOI222XL U1026 ( .A(N12814), .B(n1706), .C(n1707), .D(N12773), .E(N12805), 
        .F(n1708), .Y(n1237) );
  AOI222XL U1027 ( .A(N12811), .B(n1706), .C(n1707), .D(N12770), .E(N12802), 
        .F(n1708), .Y(n1240) );
  AOI222XL U1028 ( .A(N12813), .B(n1706), .C(n1707), .D(N12772), .E(N12804), 
        .F(n1708), .Y(n1238) );
  AOI222XL U1029 ( .A(N12810), .B(n1706), .C(n1707), .D(N12769), .E(N12801), 
        .F(n1708), .Y(n1241) );
  OAI31XL U1030 ( .A(n1885), .B(n1291), .C(cs_run), .D(n1293), .Y(n1773) );
  INVX1 U1031 ( .A(n728), .Y(n2016) );
  OAI221X1 U1032 ( .A(n1702), .B(n1131), .C(n1713), .D(n369), .E(n1723), .Y(
        n728) );
  OA222X1 U1033 ( .A(n1241), .B(n1703), .C(n2071), .D(n1705), .E(n2129), .F(
        n1704), .Y(n1723) );
  AND3X1 U1034 ( .A(n1958), .B(n1734), .C(n1957), .Y(n1670) );
  NOR2X1 U1035 ( .A(n9), .B(n449), .Y(n892) );
  XNOR2XL U1036 ( .A(n2182), .B(n2180), .Y(adder_out[5]) );
  XNOR2XL U1037 ( .A(N11546), .B(N11527), .Y(n2182) );
  XNOR2XL U1038 ( .A(N11526), .B(n2183), .Y(adder_out[4]) );
  XNOR2XL U1039 ( .A(N11555), .B(N11545), .Y(n2183) );
  OAI21X1 U1040 ( .B(n1372), .C(n2158), .A(n1373), .Y(N11527) );
  NOR2X1 U1041 ( .A(n1958), .B(instr[0]), .Y(n1167) );
  INVX1 U1042 ( .A(n739), .Y(n1423) );
  NAND3X1 U1043 ( .A(n1724), .B(n1703), .C(n2038), .Y(n1704) );
  NAND3X1 U1044 ( .A(n1575), .B(n1703), .C(n1724), .Y(n1705) );
  OAI21X1 U1045 ( .B(n1372), .C(n2156), .A(n1379), .Y(N11526) );
  NOR2X1 U1046 ( .A(n1157), .B(n429), .Y(n1611) );
  INVX1 U1047 ( .A(n449), .Y(n446) );
  NAND3X1 U1048 ( .A(n1221), .B(n1222), .C(n1929), .Y(n1185) );
  INVX1 U1049 ( .A(n375), .Y(n381) );
  INVX1 U1050 ( .A(N353), .Y(n375) );
  INVX1 U1051 ( .A(n1117), .Y(n2030) );
  INVX1 U1052 ( .A(n448), .Y(instr[5]) );
  INVX1 U1053 ( .A(n930), .Y(n2028) );
  INVX1 U1054 ( .A(n445), .Y(instr[0]) );
  INVX1 U1055 ( .A(n445), .Y(n444) );
  NOR2X1 U1056 ( .A(n1689), .B(n442), .Y(n1734) );
  ENOX1 U1057 ( .A(n671), .B(n1382), .C(n1904), .D(N12474), .Y(N11503) );
  ENOX1 U1058 ( .A(n670), .B(n1382), .C(n1904), .D(N12475), .Y(N11504) );
  AOI31X1 U1059 ( .A(n1526), .B(n196), .C(n1525), .D(n1524), .Y(n1527) );
  MUX2X1 U1060 ( .D0(n1584), .D1(n1576), .S(n175), .Y(n1525) );
  OA222X1 U1061 ( .A(n1547), .B(n1563), .C(n841), .D(n1565), .E(n2168), .F(
        n192), .Y(n165) );
  AO222X1 U1062 ( .A(N12817), .B(n1706), .C(n1707), .D(N12776), .E(N12808), 
        .F(n1708), .Y(n166) );
  INVX1 U1063 ( .A(n1812), .Y(n2122) );
  INVX1 U1064 ( .A(n1809), .Y(n2137) );
  NAND21X1 U1065 ( .B(n449), .A(n15), .Y(n2088) );
  NAND21X1 U1066 ( .B(n444), .A(n1958), .Y(n2039) );
  NAND21X1 U1067 ( .B(n1956), .A(n446), .Y(n960) );
  NOR43XL U1068 ( .B(n1357), .C(n1358), .D(n2044), .A(n1919), .Y(n1194) );
  NOR43XL U1069 ( .B(n1363), .C(n1364), .D(n1365), .A(n1366), .Y(n1357) );
  AOI21X1 U1070 ( .B(n1360), .C(n1929), .A(n1917), .Y(n1358) );
  NAND21X1 U1071 ( .B(n1808), .A(n1049), .Y(n720) );
  NAND21X1 U1072 ( .B(n1804), .A(n1047), .Y(n1049) );
  NAND21X1 U1073 ( .B(n725), .A(n1050), .Y(n1047) );
  NAND32X1 U1074 ( .B(n488), .C(n487), .A(n1654), .Y(n1176) );
  NAND21X1 U1075 ( .B(n1694), .A(n1957), .Y(n2043) );
  NAND21X1 U1076 ( .B(n2078), .A(n946), .Y(n815) );
  NAND21X1 U1077 ( .B(n1653), .A(n1929), .Y(n2044) );
  OR3XL U1078 ( .A(n528), .B(n1507), .C(n1657), .Y(n604) );
  MUX2AXL U1079 ( .D0(rn[2]), .D1(n2120), .S(n580), .Y(n865) );
  MUX2X1 U1080 ( .D0(n318), .D1(n313), .S(n2066), .Y(rn[2]) );
  MUX4X1 U1081 ( .D0(n317), .D1(n315), .D2(n316), .D3(n314), .S0(n114), .S1(
        n101), .Y(n318) );
  MUX4X1 U1082 ( .D0(n312), .D1(n310), .D2(n311), .D3(n309), .S0(n114), .S1(
        n101), .Y(n313) );
  OR3XL U1083 ( .A(n527), .B(n191), .C(n1360), .Y(n1507) );
  INVX1 U1084 ( .A(n1189), .Y(n2065) );
  NAND31X1 U1085 ( .C(n1507), .A(n1658), .B(n1657), .Y(n1508) );
  INVX1 U1086 ( .A(n1050), .Y(n1274) );
  NOR21XL U1087 ( .B(n1713), .A(n1725), .Y(n1724) );
  AOI222XL U1088 ( .A(N12815), .B(n1706), .C(n1707), .D(N12774), .E(N12806), 
        .F(n1708), .Y(n1236) );
  AOI222XL U1089 ( .A(N12816), .B(n1706), .C(n1707), .D(N12775), .E(N12807), 
        .F(n1708), .Y(n1235) );
  AOI222XL U1090 ( .A(N12812), .B(n1706), .C(n1707), .D(N12771), .E(N12803), 
        .F(n1708), .Y(n1239) );
  INVX1 U1091 ( .A(n1718), .Y(n1989) );
  OAI221X1 U1092 ( .A(n865), .B(n1702), .C(n1713), .D(n64), .E(n1719), .Y(
        n1718) );
  OA222X1 U1093 ( .A(n1239), .B(n1703), .C(n2121), .D(n1705), .E(n1964), .F(
        n1704), .Y(n1719) );
  NAND21X1 U1094 ( .B(n1654), .A(n1927), .Y(n1186) );
  INVX1 U1095 ( .A(n1188), .Y(n2066) );
  NAND41X1 U1096 ( .D(n1658), .A(n1929), .B(n1928), .C(n1657), .Y(n1179) );
  INVX1 U1097 ( .A(n1507), .Y(n1928) );
  NAND3X1 U1098 ( .A(n1731), .B(n1957), .C(intcall), .Y(n1499) );
  NAND4X1 U1099 ( .A(n1650), .B(n1647), .C(n1651), .D(n1652), .Y(n1365) );
  NOR2X1 U1100 ( .A(n1955), .B(n446), .Y(n1119) );
  INVX1 U1101 ( .A(n433), .Y(n429) );
  INVX1 U1102 ( .A(n2077), .Y(n433) );
  INVX1 U1103 ( .A(n1821), .Y(n2080) );
  AND2X1 U1104 ( .A(n401), .B(n1474), .Y(N582) );
  NOR2X1 U1105 ( .A(n2082), .B(n2105), .Y(n1594) );
  INVX1 U1106 ( .A(n509), .Y(n1944) );
  INVX1 U1107 ( .A(ramdatai[0]), .Y(n648) );
  INVX1 U1108 ( .A(n1124), .Y(n2100) );
  INVX1 U1109 ( .A(n1566), .Y(n2010) );
  INVX1 U1110 ( .A(n1509), .Y(n1221) );
  NAND32X1 U1111 ( .B(n1735), .C(n1508), .A(n1654), .Y(n1509) );
  INVX1 U1112 ( .A(n440), .Y(dps[1]) );
  INVX1 U1113 ( .A(ramdatai[1]), .Y(n2173) );
  NOR2X1 U1114 ( .A(n2105), .B(n1955), .Y(n1593) );
  NOR4XL U1115 ( .A(n1215), .B(n1216), .C(n1217), .D(n1201), .Y(n1203) );
  NAND41X1 U1116 ( .D(n1918), .A(n1226), .B(n1186), .C(n1227), .Y(n1215) );
  OAI21X1 U1117 ( .B(n1218), .C(n1219), .A(n1194), .Y(n1216) );
  INVX1 U1118 ( .A(n1666), .Y(n1918) );
  INVX1 U1119 ( .A(n370), .Y(n369) );
  ENOX1 U1120 ( .A(n672), .B(n1382), .C(n1904), .D(N12473), .Y(N11502) );
  INVX1 U1121 ( .A(n901), .Y(n2097) );
  NAND3X1 U1122 ( .A(n1167), .B(n2106), .C(n1922), .Y(n1694) );
  NAND2X1 U1123 ( .A(n452), .B(n683), .Y(n681) );
  OAI21X1 U1124 ( .B(n1885), .C(n684), .A(n680), .Y(n683) );
  INVX1 U1125 ( .A(n1224), .Y(n521) );
  INVX1 U1126 ( .A(n1226), .Y(n529) );
  INVX1 U1127 ( .A(n1653), .Y(n527) );
  NOR32XL U1128 ( .B(n1647), .C(n1648), .A(n1649), .Y(n1366) );
  NOR21XL U1129 ( .B(n1740), .A(n2092), .Y(n908) );
  NAND31X1 U1130 ( .C(n1005), .A(n1943), .B(n1010), .Y(n1032) );
  NAND21X1 U1131 ( .B(n2100), .A(n1839), .Y(n1159) );
  NAND32X1 U1132 ( .B(n1956), .C(n2037), .A(n1946), .Y(n2035) );
  OR2X1 U1133 ( .A(n125), .B(n167), .Y(n629) );
  AOI21X1 U1134 ( .B(n1910), .C(n15), .A(n1344), .Y(n167) );
  NOR32XL U1135 ( .B(n1220), .C(n2046), .A(n1228), .Y(n1217) );
  NAND32X1 U1136 ( .B(n528), .C(n527), .A(n191), .Y(n560) );
  NAND21X1 U1137 ( .B(n2093), .A(n576), .Y(n1581) );
  NAND21X1 U1138 ( .B(n1006), .A(n1942), .Y(n686) );
  NAND21X1 U1139 ( .B(n2093), .A(n1017), .Y(n1582) );
  OAI21X1 U1140 ( .B(n1372), .C(n2139), .A(n1373), .Y(N11528) );
  NOR3XL U1141 ( .A(n2042), .B(n2100), .C(n1821), .Y(n168) );
  XNOR3X1 U1142 ( .A(N11541), .B(N11549), .C(N11522), .Y(n544) );
  OAI22X1 U1143 ( .A(n1579), .B(n2078), .C(n430), .D(n1580), .Y(n646) );
  AND2X1 U1144 ( .A(n1734), .B(n903), .Y(n1062) );
  OAI32X1 U1145 ( .A(n2101), .B(n1736), .C(n123), .D(n430), .E(n1600), .Y(
        n1725) );
  OA22X1 U1146 ( .A(n2127), .B(n1183), .C(n1176), .D(n2159), .Y(n605) );
  OA22X1 U1147 ( .A(n1183), .B(n783), .C(n1176), .D(n2140), .Y(n558) );
  XNOR3X1 U1148 ( .A(N11523), .B(N11542), .C(n530), .Y(n531) );
  NOR2X1 U1149 ( .A(n442), .B(n1958), .Y(n1599) );
  NOR2X1 U1150 ( .A(n2106), .B(n1956), .Y(n1116) );
  NOR2X1 U1151 ( .A(n2104), .B(n123), .Y(intcall) );
  NOR2X1 U1152 ( .A(n2101), .B(n2106), .Y(n1489) );
  NOR2X1 U1153 ( .A(n2105), .B(n2100), .Y(n1331) );
  NAND2X1 U1154 ( .A(n1713), .B(n1725), .Y(n1702) );
  NOR2X1 U1155 ( .A(n2098), .B(n448), .Y(n1597) );
  INVX1 U1156 ( .A(n1941), .Y(n2072) );
  INVX1 U1157 ( .A(n369), .Y(n374) );
  NOR42XL U1158 ( .C(n1209), .D(n1220), .A(n1185), .B(n1211), .Y(n1201) );
  NOR2X1 U1159 ( .A(n737), .B(n370), .Y(n1673) );
  INVX1 U1160 ( .A(n1804), .Y(codefetch_s) );
  INVX1 U1161 ( .A(n626), .Y(n1565) );
  NAND21X1 U1162 ( .B(n194), .A(n629), .Y(n626) );
  NOR3XL U1163 ( .A(n2049), .B(n2050), .C(n1650), .Y(n1648) );
  INVX1 U1164 ( .A(n2081), .Y(n1605) );
  AND2X1 U1165 ( .A(n391), .B(n1401), .Y(N11501) );
  NAND3X1 U1166 ( .A(n912), .B(n1117), .C(n2080), .Y(n972) );
  INVX1 U1167 ( .A(n570), .Y(n1017) );
  NAND21X1 U1168 ( .B(n449), .A(n1673), .Y(n570) );
  INVX1 U1169 ( .A(n487), .Y(n1735) );
  NAND2X1 U1170 ( .A(n1609), .B(n10), .Y(n1680) );
  INVX1 U1171 ( .A(n2077), .Y(n432) );
  INVX1 U1172 ( .A(n903), .Y(n2101) );
  ENOX1 U1173 ( .A(n673), .B(n1382), .C(n1904), .D(N12471), .Y(N11500) );
  NAND2X1 U1174 ( .A(n1835), .B(n1946), .Y(n1608) );
  NAND2X1 U1175 ( .A(n1598), .B(n1062), .Y(n1579) );
  OA22X1 U1176 ( .A(n2078), .B(n1585), .C(n431), .D(n1586), .Y(n169) );
  OA22X1 U1177 ( .A(n2078), .B(n1577), .C(n431), .D(n1578), .Y(n170) );
  INVX1 U1178 ( .A(n1652), .Y(n2050) );
  INVX1 U1179 ( .A(n1651), .Y(n2049) );
  NAND21X1 U1180 ( .B(n624), .A(n194), .Y(n1422) );
  NAND43X1 U1181 ( .B(n1422), .C(n643), .D(n707), .A(n642), .Y(n1539) );
  OR4X1 U1182 ( .A(n1424), .B(n1422), .C(n707), .D(n171), .Y(n1515) );
  NAND4X1 U1183 ( .A(n1457), .B(n1553), .C(n1540), .D(n1458), .Y(n171) );
  NAND21X1 U1184 ( .B(n1660), .A(n1920), .Y(n1666) );
  OR2X1 U1185 ( .A(n2078), .B(n1158), .Y(n618) );
  NAND5XL U1186 ( .A(n644), .B(n1537), .C(n643), .D(n1456), .E(n642), .Y(n1553) );
  OAI21BBX1 U1187 ( .A(n1916), .B(n1961), .C(n1470), .Y(n1494) );
  NAND21X1 U1188 ( .B(n2093), .A(n1599), .Y(n612) );
  NAND32X1 U1189 ( .B(n538), .C(n537), .A(n536), .Y(n1511) );
  NAND21X1 U1190 ( .B(n1961), .A(n1916), .Y(n1510) );
  NAND21X1 U1191 ( .B(n2093), .A(n1948), .Y(n601) );
  NAND32X1 U1192 ( .B(n524), .C(n523), .A(n522), .Y(n541) );
  INVX1 U1193 ( .A(n1223), .Y(n522) );
  INVX1 U1194 ( .A(n1660), .Y(n523) );
  INVX1 U1195 ( .A(n520), .Y(n1916) );
  NAND21X1 U1196 ( .B(n1618), .A(n552), .Y(n520) );
  NAND21X1 U1197 ( .B(n1961), .A(n630), .Y(n1563) );
  AOI222XL U1198 ( .A(n369), .B(n1593), .C(n2105), .D(n1689), .E(n2104), .F(
        n10), .Y(n1858) );
  NAND32X1 U1199 ( .B(n518), .C(n538), .A(n536), .Y(n1467) );
  INVX1 U1200 ( .A(n537), .Y(n518) );
  NAND42X1 U1201 ( .C(n1211), .D(n1213), .A(n1220), .B(n1221), .Y(n1219) );
  XNOR2XL U1202 ( .A(n1370), .B(n1966), .Y(n1230) );
  NAND32X1 U1203 ( .B(n1387), .C(n514), .A(n513), .Y(n538) );
  INVX1 U1204 ( .A(n1614), .Y(n513) );
  INVX1 U1205 ( .A(n1618), .Y(n514) );
  OAI221X1 U1206 ( .A(n16), .B(n633), .C(n431), .D(n4), .E(n1552), .Y(n756) );
  OA22X1 U1207 ( .A(n124), .B(n632), .C(n430), .D(n631), .Y(n633) );
  INVX1 U1208 ( .A(n1609), .Y(n631) );
  NAND2X1 U1209 ( .A(n370), .B(n1860), .Y(n916) );
  INVX1 U1210 ( .A(n1569), .Y(n1552) );
  NAND2X1 U1211 ( .A(n1014), .B(n1942), .Y(n1275) );
  NOR3XL U1212 ( .A(n2097), .B(n1958), .C(n2092), .Y(n1674) );
  OAI32X1 U1213 ( .A(n916), .B(n1858), .C(n449), .D(n1859), .E(n1955), .Y(
        n1856) );
  AOI32X1 U1214 ( .A(n2020), .B(n1958), .C(n912), .D(n1686), .E(n1857), .Y(
        n1859) );
  INVX1 U1215 ( .A(n1858), .Y(n2020) );
  INVX1 U1216 ( .A(n1387), .Y(n552) );
  INVX1 U1217 ( .A(n1303), .Y(n1526) );
  INVX1 U1218 ( .A(n2019), .Y(n1940) );
  OAI31XL U1219 ( .A(n2102), .B(n10), .C(n2030), .D(n2029), .Y(n1751) );
  INVX1 U1220 ( .A(n1835), .Y(n2029) );
  NOR2X1 U1221 ( .A(n1061), .B(n1839), .Y(n1112) );
  AND2XL U1222 ( .A(n400), .B(n1301), .Y(N11499) );
  NOR21XL U1223 ( .B(n1822), .A(n2088), .Y(n1793) );
  NAND21X1 U1224 ( .B(n1957), .A(n950), .Y(n2096) );
  NAND21X1 U1225 ( .B(n21), .A(n739), .Y(n635) );
  NAND21X1 U1226 ( .B(n1387), .A(n1614), .Y(n1512) );
  NAND31X1 U1227 ( .C(n1303), .A(n663), .B(n1411), .Y(n664) );
  MUX2IX1 U1228 ( .D0(n660), .D1(n659), .S(n657), .Y(n663) );
  INVX1 U1229 ( .A(n1576), .Y(n659) );
  INVX1 U1230 ( .A(n1584), .Y(n660) );
  NAND21X1 U1231 ( .B(n1957), .A(n1911), .Y(n632) );
  AOI211X1 U1232 ( .C(n1619), .D(n1620), .A(n89), .B(n125), .Y(n1614) );
  AOI211X1 U1233 ( .C(n1956), .D(n891), .A(n1598), .B(n1061), .Y(n1620) );
  NOR3XL U1234 ( .A(n2080), .B(n1952), .C(n1922), .Y(n1619) );
  MUX2AXL U1235 ( .D0(n2163), .D1(n1453), .S(n450), .Y(ramsfraddr_comb[4]) );
  OAI31XL U1236 ( .A(n612), .B(n124), .C(n999), .D(n615), .Y(n603) );
  AND2X1 U1237 ( .A(n1860), .B(n442), .Y(n1834) );
  INVX1 U1238 ( .A(n615), .Y(n622) );
  AND4X1 U1239 ( .A(n904), .B(n905), .C(n906), .D(n907), .Y(n884) );
  AOI211X1 U1240 ( .C(n912), .D(n913), .A(n914), .B(n915), .Y(n906) );
  NOR4XL U1241 ( .A(n908), .B(n909), .C(n910), .D(n911), .Y(n907) );
  NOR3XL U1242 ( .A(n922), .B(n923), .C(n924), .Y(n904) );
  XNOR2XL U1243 ( .A(n1057), .B(n1970), .Y(n1053) );
  XNOR2XL U1244 ( .A(n1055), .B(n1056), .Y(n1054) );
  INVX1 U1245 ( .A(n634), .Y(n1571) );
  NAND21X1 U1246 ( .B(n2078), .A(n924), .Y(n634) );
  NOR3XL U1247 ( .A(n16), .B(n1911), .C(n2037), .Y(n1162) );
  AND2X1 U1248 ( .A(n1061), .B(n1835), .Y(n1787) );
  NOR2X1 U1249 ( .A(n2105), .B(n446), .Y(n1631) );
  OAI21X1 U1250 ( .B(n1372), .C(n2160), .A(n1379), .Y(n1232) );
  INVX1 U1251 ( .A(n793), .Y(n772) );
  OAI31XL U1252 ( .A(n2039), .B(n125), .C(n809), .D(n1244), .Y(n1634) );
  OAI21X1 U1253 ( .B(n2092), .C(n896), .A(n2091), .Y(n1152) );
  OAI21X1 U1254 ( .B(n2083), .C(n896), .A(n1639), .Y(n1625) );
  AND2X1 U1255 ( .A(n392), .B(n557), .Y(N12905) );
  XOR3X1 U1256 ( .A(n1048), .B(n1051), .C(n556), .Y(n557) );
  XNOR2XL U1257 ( .A(n1994), .B(n1893), .Y(n1051) );
  XNOR2XL U1258 ( .A(n1053), .B(n1054), .Y(n1048) );
  NOR2X1 U1259 ( .A(n1956), .B(n1957), .Y(n1118) );
  MUX2IX1 U1260 ( .D0(n2127), .D1(n2151), .S(n1571), .Y(n172) );
  INVX1 U1261 ( .A(n912), .Y(n2102) );
  OAI21X1 U1262 ( .B(n1114), .C(n64), .A(n1115), .Y(n1626) );
  INVX1 U1263 ( .A(n1026), .Y(n777) );
  NAND21X1 U1264 ( .B(n2099), .A(n1332), .Y(n1244) );
  OAI32X1 U1265 ( .A(n2033), .B(n2068), .C(n1954), .D(n1333), .E(n2077), .Y(
        n1332) );
  AOI32X1 U1266 ( .A(n891), .B(n120), .C(n1948), .D(n1899), .E(n2068), .Y(
        n1333) );
  INVX1 U1267 ( .A(n2033), .Y(n1899) );
  AOI22AXL U1268 ( .A(n1123), .B(n2190), .D(n1114), .C(n901), .Y(n1629) );
  NAND2X1 U1269 ( .A(n1910), .B(n1682), .Y(n1638) );
  INVX1 U1270 ( .A(n736), .Y(n2068) );
  NOR3XL U1271 ( .A(n2039), .B(n16), .C(n1858), .Y(n1861) );
  NAND2X1 U1272 ( .A(n1214), .B(n1228), .Y(n1211) );
  OAI211X1 U1273 ( .C(n1594), .D(n1946), .A(n1117), .B(n912), .Y(n1679) );
  INVX1 U1274 ( .A(n902), .Y(n2083) );
  NAND2X1 U1275 ( .A(n1598), .B(n2041), .Y(n1781) );
  AOI31X1 U1276 ( .A(n884), .B(n885), .C(n2031), .D(n124), .Y(n883) );
  INVX1 U1277 ( .A(n886), .Y(n2031) );
  NAND2X1 U1278 ( .A(n1822), .B(n1598), .Y(n1776) );
  NAND2X1 U1279 ( .A(n1598), .B(n1835), .Y(n1777) );
  NAND2X1 U1280 ( .A(n1834), .B(n902), .Y(n1771) );
  NAND2X1 U1281 ( .A(n446), .B(n57), .Y(n1114) );
  INVX1 U1282 ( .A(n1297), .Y(n2017) );
  NAND4X1 U1283 ( .A(n1212), .B(n1222), .C(n1223), .D(n1224), .Y(n1218) );
  NAND2X1 U1284 ( .A(n1740), .B(n1682), .Y(n1752) );
  NAND2X1 U1285 ( .A(n1892), .B(n1839), .Y(n1639) );
  NAND2X1 U1286 ( .A(n884), .B(n899), .Y(n749) );
  OAI31XL U1287 ( .A(n900), .B(n901), .C(n902), .D(n903), .Y(n899) );
  OAI22X1 U1288 ( .A(instr[5]), .B(n2095), .C(n16), .D(n64), .Y(n900) );
  INVX1 U1289 ( .A(n1684), .Y(n1893) );
  NAND2X1 U1290 ( .A(n1599), .B(n2106), .Y(n1871) );
  OR2X1 U1291 ( .A(n737), .B(n2083), .Y(n1755) );
  NOR21XL U1292 ( .B(n1206), .A(n1207), .Y(n1220) );
  NAND32X1 U1293 ( .B(n430), .C(n517), .A(n516), .Y(n536) );
  INVX1 U1294 ( .A(n1489), .Y(n517) );
  OAI221X1 U1295 ( .A(n1956), .B(n515), .C(n63), .D(n950), .E(n2088), .Y(n516)
         );
  INVX1 U1296 ( .A(n1631), .Y(n515) );
  NAND43X1 U1297 ( .B(n635), .C(n582), .D(n1909), .A(n636), .Y(n1457) );
  INVX1 U1298 ( .A(n1602), .Y(n582) );
  NAND32X1 U1299 ( .B(n63), .C(n2039), .A(n950), .Y(n2033) );
  MUX2X1 U1300 ( .D0(n783), .D1(n2129), .S(n1571), .Y(n656) );
  NAND21X1 U1301 ( .B(n2093), .A(n1021), .Y(n1760) );
  NAND21X1 U1302 ( .B(n1026), .A(n1022), .Y(n1758) );
  INVX1 U1303 ( .A(n936), .Y(N12473) );
  NAND21X1 U1304 ( .B(n1808), .A(n1056), .Y(n936) );
  NOR21XL U1305 ( .B(n1822), .A(n2092), .Y(n1788) );
  NAND21X1 U1306 ( .B(n1457), .A(pc_i[0]), .Y(n641) );
  AND2X1 U1307 ( .A(n1599), .B(n1124), .Y(n1828) );
  INVX1 U1308 ( .A(pc_i[9]), .Y(n984) );
  NAND21X1 U1309 ( .B(n1908), .A(n784), .Y(n1421) );
  MUX2AXL U1310 ( .D0(n2132), .D1(n1452), .S(n450), .Y(ramsfraddr_comb[3]) );
  NAND21X1 U1311 ( .B(n782), .A(n1757), .Y(n792) );
  NOR2X1 U1312 ( .A(n930), .B(n22), .Y(n1424) );
  AND2X1 U1313 ( .A(n1834), .B(n1598), .Y(n1782) );
  AND2X1 U1314 ( .A(n1822), .B(n1061), .Y(n1786) );
  OAI211X1 U1315 ( .C(n2095), .D(n1875), .A(n972), .B(n2091), .Y(n1163) );
  NAND2X1 U1316 ( .A(n892), .B(n69), .Y(n1875) );
  INVX1 U1317 ( .A(n2098), .Y(n1895) );
  INVX1 U1318 ( .A(n637), .Y(n642) );
  NAND21X1 U1319 ( .B(n1602), .A(n636), .Y(n637) );
  NAND42X1 U1320 ( .C(n918), .D(n1845), .A(n1846), .B(n717), .Y(n1844) );
  AOI22X1 U1321 ( .A(n1489), .B(n960), .C(n1848), .D(n89), .Y(n1846) );
  NAND41X1 U1322 ( .D(n915), .A(n1752), .B(n1755), .C(n1851), .Y(n1845) );
  OAI222XL U1323 ( .A(n1849), .B(n2030), .C(n1850), .D(n2106), .E(instr[5]), 
        .F(n1115), .Y(n1848) );
  AOI21X1 U1324 ( .B(n1839), .C(n369), .A(n1922), .Y(n1850) );
  AOI31X1 U1325 ( .A(n1922), .B(n442), .C(n1124), .D(n1163), .Y(n1874) );
  OAI211X1 U1326 ( .C(n797), .D(n796), .A(n794), .B(n949), .Y(n798) );
  AND3X1 U1327 ( .A(n1026), .B(n999), .C(n793), .Y(n797) );
  INVX1 U1328 ( .A(n993), .Y(n1888) );
  NAND21X1 U1329 ( .B(n2093), .A(n992), .Y(n993) );
  NAND3X1 U1330 ( .A(n89), .B(n1956), .C(n932), .Y(n1125) );
  NAND3X1 U1331 ( .A(n1125), .B(n1157), .C(n1158), .Y(n919) );
  INVX1 U1332 ( .A(n851), .Y(N12474) );
  NAND21X1 U1333 ( .B(n398), .A(n1055), .Y(n851) );
  INVX1 U1334 ( .A(n565), .Y(N12471) );
  NAND21X1 U1335 ( .B(n1994), .A(n387), .Y(n565) );
  INVX1 U1336 ( .A(n567), .Y(N12476) );
  NAND21X1 U1337 ( .B(n1970), .A(n388), .Y(n567) );
  NAND3X1 U1338 ( .A(n1948), .B(n64), .C(n2080), .Y(n1693) );
  INVX1 U1339 ( .A(n1667), .Y(n2018) );
  NAND32X1 U1340 ( .B(n16), .C(n2037), .A(n950), .Y(n791) );
  INVX1 U1341 ( .A(n483), .Y(n1460) );
  NAND21X1 U1342 ( .B(n125), .A(n1938), .Y(n483) );
  INVX1 U1343 ( .A(n937), .Y(N12475) );
  NAND21X1 U1344 ( .B(n1808), .A(n1057), .Y(n937) );
  OAI211X1 U1345 ( .C(n2039), .D(n1159), .A(n949), .B(n2081), .Y(n886) );
  NAND21X1 U1346 ( .B(n1908), .A(n786), .Y(n1411) );
  AND2X1 U1347 ( .A(n391), .B(n1684), .Y(N12472) );
  INVX1 U1348 ( .A(n506), .Y(n1938) );
  INVX1 U1349 ( .A(n1757), .Y(n911) );
  NAND2X1 U1350 ( .A(n1834), .B(n10), .Y(n897) );
  NAND21X1 U1351 ( .B(n2141), .A(n388), .Y(n2002) );
  NAND21X1 U1352 ( .B(n2128), .A(n388), .Y(n2004) );
  NAND21X1 U1353 ( .B(n2134), .A(n388), .Y(n2003) );
  NAND21X1 U1354 ( .B(n2120), .A(n387), .Y(n2005) );
  NAND21X1 U1355 ( .B(n1610), .A(n849), .Y(n973) );
  NAND21X1 U1356 ( .B(n795), .A(n849), .Y(n974) );
  NAND32X1 U1357 ( .B(n1896), .C(n834), .A(n833), .Y(n843) );
  NAND21X1 U1358 ( .B(n2064), .A(n387), .Y(n2006) );
  NAND21X1 U1359 ( .B(n2136), .A(n388), .Y(n2001) );
  NAND21X1 U1360 ( .B(n2053), .A(n387), .Y(n2007) );
  INVX1 U1361 ( .A(n784), .Y(n1433) );
  INVX1 U1362 ( .A(n786), .Y(n1415) );
  INVX1 U1363 ( .A(n1606), .Y(n1529) );
  OAI22XL U1364 ( .A(n459), .B(n827), .C(n1130), .D(n1564), .Y(N12721) );
  AOI221XL U1365 ( .A(n970), .B(n962), .C(n1132), .D(ramdatai[7]), .E(n1133), 
        .Y(n827) );
  OAI22X1 U1366 ( .A(n2021), .B(n1999), .C(n17), .D(n1134), .Y(n1133) );
  OAI22XL U1367 ( .A(n459), .B(n966), .C(n1130), .D(n965), .Y(N12714) );
  AOI221XL U1368 ( .A(n963), .B(n962), .C(n1132), .D(ramdatai[0]), .E(n1150), 
        .Y(n966) );
  OAI22X1 U1369 ( .A(n2021), .B(n1991), .C(n31), .D(n1134), .Y(n1150) );
  NAND21X1 U1370 ( .B(n124), .A(n915), .Y(n837) );
  NAND21X1 U1371 ( .B(n2130), .A(n388), .Y(n2000) );
  NAND32X1 U1372 ( .B(n398), .C(finishdiv), .A(n467), .Y(n486) );
  INVX1 U1373 ( .A(n1222), .Y(n467) );
  INVX1 U1374 ( .A(n810), .Y(n1897) );
  NAND32X1 U1375 ( .B(n125), .C(n69), .A(n1945), .Y(n810) );
  NAND2X1 U1376 ( .A(n933), .B(n932), .Y(n833) );
  INVX1 U1377 ( .A(pc_i[1]), .Y(n987) );
  INVX1 U1378 ( .A(n602), .Y(n1894) );
  NAND21X1 U1379 ( .B(n2161), .A(n808), .Y(n602) );
  NAND21X1 U1380 ( .B(n1804), .A(n387), .Y(n722) );
  AO21X1 U1381 ( .B(n395), .C(n476), .A(n462), .Y(N11491) );
  INVX1 U1382 ( .A(n1662), .Y(n476) );
  INVX1 U1383 ( .A(n1664), .Y(n1246) );
  NAND43X1 U1384 ( .B(n1663), .C(n396), .D(n1661), .A(n1012), .Y(n1664) );
  INVX1 U1385 ( .A(n1015), .Y(n1661) );
  AND2X1 U1386 ( .A(N10579), .B(n2019), .Y(N371) );
  AND2X1 U1387 ( .A(N10580), .B(n2019), .Y(N372) );
  INVX1 U1388 ( .A(n1722), .Y(n1007) );
  NAND21X1 U1389 ( .B(n8), .A(n388), .Y(n1722) );
  NAND2X1 U1390 ( .A(n1007), .B(n1012), .Y(n1011) );
  NAND2X1 U1391 ( .A(n1007), .B(n1010), .Y(n1009) );
  OAI221X1 U1392 ( .A(n2150), .B(n1342), .C(n795), .D(n2007), .E(n457), .Y(
        N12485) );
  OAI221X1 U1393 ( .A(n2149), .B(n1342), .C(n2006), .D(n795), .E(n457), .Y(
        N12486) );
  OAI221X1 U1394 ( .A(n2148), .B(n1342), .C(n2005), .D(n795), .E(n456), .Y(
        N12487) );
  OAI22X1 U1395 ( .A(n926), .B(n85), .C(n2032), .D(n1256), .Y(N12602) );
  OAI22X1 U1396 ( .A(n848), .B(n85), .C(n1984), .D(n97), .Y(N12607) );
  OAI22X1 U1397 ( .A(n807), .B(n85), .C(n1979), .D(n97), .Y(N12532) );
  OAI22X1 U1398 ( .A(n801), .B(n85), .C(n1978), .D(n97), .Y(N12533) );
  OAI22X1 U1399 ( .A(n790), .B(n85), .C(n1977), .D(n97), .Y(N12534) );
  OAI22X1 U1400 ( .A(n785), .B(n85), .C(n1976), .D(n97), .Y(N12535) );
  OAI22X1 U1401 ( .A(n780), .B(n85), .C(n1975), .D(n97), .Y(N12536) );
  OAI22X1 U1402 ( .A(n775), .B(n85), .C(n1974), .D(n97), .Y(N12537) );
  OAI22X1 U1403 ( .A(n926), .B(n96), .C(n2032), .D(n1254), .Y(N12611) );
  OAI22X1 U1404 ( .A(n848), .B(n96), .C(n1984), .D(n83), .Y(N12616) );
  OAI22X1 U1405 ( .A(n807), .B(n96), .C(n1979), .D(n83), .Y(N12541) );
  OAI22X1 U1406 ( .A(n801), .B(n96), .C(n1978), .D(n83), .Y(N12542) );
  OAI22X1 U1407 ( .A(n790), .B(n96), .C(n1977), .D(n83), .Y(N12543) );
  OAI22X1 U1408 ( .A(n785), .B(n96), .C(n1976), .D(n83), .Y(N12544) );
  OAI22X1 U1409 ( .A(n780), .B(n96), .C(n1975), .D(n83), .Y(N12545) );
  OAI22X1 U1410 ( .A(n775), .B(n96), .C(n1974), .D(n83), .Y(N12546) );
  OAI22X1 U1411 ( .A(n926), .B(n68), .C(n2032), .D(n1252), .Y(N12620) );
  OAI22X1 U1412 ( .A(n848), .B(n68), .C(n1984), .D(n76), .Y(N12625) );
  OAI22X1 U1413 ( .A(n807), .B(n68), .C(n1979), .D(n76), .Y(N12550) );
  OAI22X1 U1414 ( .A(n801), .B(n68), .C(n1978), .D(n76), .Y(N12551) );
  OAI22X1 U1415 ( .A(n790), .B(n68), .C(n1977), .D(n76), .Y(N12552) );
  OAI22X1 U1416 ( .A(n785), .B(n68), .C(n1976), .D(n76), .Y(N12553) );
  OAI22X1 U1417 ( .A(n780), .B(n68), .C(n1975), .D(n76), .Y(N12554) );
  OAI22X1 U1418 ( .A(n775), .B(n68), .C(n1974), .D(n76), .Y(N12555) );
  OAI22X1 U1419 ( .A(n926), .B(n75), .C(n2032), .D(n1250), .Y(N12629) );
  OAI22X1 U1420 ( .A(n848), .B(n75), .C(n1984), .D(n66), .Y(N12634) );
  OAI22X1 U1421 ( .A(n807), .B(n75), .C(n1979), .D(n66), .Y(N12559) );
  OAI22X1 U1422 ( .A(n801), .B(n75), .C(n1978), .D(n66), .Y(N12560) );
  OAI22X1 U1423 ( .A(n790), .B(n75), .C(n1977), .D(n66), .Y(N12561) );
  OAI22X1 U1424 ( .A(n785), .B(n75), .C(n1976), .D(n66), .Y(N12562) );
  OAI22X1 U1425 ( .A(n780), .B(n75), .C(n1975), .D(n66), .Y(N12563) );
  OAI22X1 U1426 ( .A(n775), .B(n75), .C(n1974), .D(n66), .Y(N12564) );
  OAI22X1 U1427 ( .A(n926), .B(n94), .C(n2032), .D(n1264), .Y(N12566) );
  OAI22X1 U1428 ( .A(n848), .B(n94), .C(n1984), .D(n110), .Y(N12571) );
  OAI22X1 U1429 ( .A(n807), .B(n94), .C(n1979), .D(n110), .Y(N12496) );
  OAI22X1 U1430 ( .A(n801), .B(n94), .C(n1978), .D(n110), .Y(N12497) );
  OAI22X1 U1431 ( .A(n790), .B(n94), .C(n1977), .D(n110), .Y(N12498) );
  OAI22X1 U1432 ( .A(n785), .B(n94), .C(n1976), .D(n110), .Y(N12499) );
  OAI22X1 U1433 ( .A(n780), .B(n94), .C(n1975), .D(n110), .Y(N12500) );
  OAI22X1 U1434 ( .A(n775), .B(n94), .C(n1974), .D(n110), .Y(N12501) );
  OAI22X1 U1435 ( .A(n926), .B(n109), .C(n2032), .D(n1262), .Y(N12575) );
  OAI22X1 U1436 ( .A(n848), .B(n109), .C(n1984), .D(n62), .Y(N12580) );
  OAI22X1 U1437 ( .A(n807), .B(n109), .C(n1979), .D(n62), .Y(N12505) );
  OAI22X1 U1438 ( .A(n801), .B(n109), .C(n1978), .D(n62), .Y(N12506) );
  OAI22X1 U1439 ( .A(n790), .B(n109), .C(n1977), .D(n62), .Y(N12507) );
  OAI22X1 U1440 ( .A(n785), .B(n109), .C(n1976), .D(n62), .Y(N12508) );
  OAI22X1 U1441 ( .A(n780), .B(n109), .C(n1975), .D(n62), .Y(N12509) );
  OAI22X1 U1442 ( .A(n775), .B(n109), .C(n1974), .D(n62), .Y(N12510) );
  OAI22X1 U1443 ( .A(n926), .B(n82), .C(n2032), .D(n1260), .Y(N12584) );
  OAI22X1 U1444 ( .A(n848), .B(n82), .C(n1984), .D(n60), .Y(N12589) );
  OAI22X1 U1445 ( .A(n807), .B(n82), .C(n1979), .D(n60), .Y(N12514) );
  OAI22X1 U1446 ( .A(n801), .B(n82), .C(n1978), .D(n60), .Y(N12515) );
  OAI22X1 U1447 ( .A(n790), .B(n82), .C(n1977), .D(n60), .Y(N12516) );
  OAI22X1 U1448 ( .A(n785), .B(n82), .C(n1976), .D(n60), .Y(N12517) );
  OAI22X1 U1449 ( .A(n780), .B(n82), .C(n1975), .D(n60), .Y(N12518) );
  OAI22X1 U1450 ( .A(n775), .B(n82), .C(n1974), .D(n60), .Y(N12519) );
  OAI22X1 U1451 ( .A(n926), .B(n73), .C(n2032), .D(n1258), .Y(N12593) );
  OAI22X1 U1452 ( .A(n848), .B(n73), .C(n1984), .D(n58), .Y(N12598) );
  OAI22X1 U1453 ( .A(n807), .B(n73), .C(n1979), .D(n58), .Y(N12523) );
  OAI22X1 U1454 ( .A(n801), .B(n73), .C(n1978), .D(n58), .Y(N12524) );
  OAI22X1 U1455 ( .A(n790), .B(n73), .C(n1977), .D(n58), .Y(N12525) );
  OAI22X1 U1456 ( .A(n785), .B(n73), .C(n1976), .D(n58), .Y(N12526) );
  OAI22X1 U1457 ( .A(n780), .B(n73), .C(n1975), .D(n58), .Y(N12527) );
  OAI22X1 U1458 ( .A(n775), .B(n73), .C(n1974), .D(n58), .Y(N12528) );
  OAI22AX1 U1459 ( .D(n1296), .C(n399), .A(n1455), .B(n997), .Y(N11487) );
  OAI21X1 U1460 ( .B(n1002), .C(n1001), .A(n453), .Y(N13284) );
  OAI21X1 U1461 ( .B(n1001), .C(n1003), .A(n453), .Y(N13257) );
  OAI21X1 U1462 ( .B(n1001), .C(n1004), .A(n453), .Y(N13248) );
  OAI21X1 U1463 ( .B(n1005), .C(n1001), .A(n454), .Y(N13239) );
  OAI21X1 U1464 ( .B(n1006), .C(n1001), .A(n453), .Y(N13230) );
  OAI21X1 U1465 ( .B(n1002), .C(n1009), .A(n453), .Y(N13212) );
  OAI21X1 U1466 ( .B(n1003), .C(n1009), .A(n454), .Y(N13185) );
  OAI21X1 U1467 ( .B(n1004), .C(n1009), .A(n454), .Y(N13176) );
  OAI21X1 U1468 ( .B(n1005), .C(n1009), .A(n454), .Y(N13167) );
  OAI21X1 U1469 ( .B(n1006), .C(n1009), .A(n454), .Y(N13158) );
  OAI21X1 U1470 ( .B(n1002), .C(n1011), .A(n454), .Y(N13140) );
  OAI21X1 U1471 ( .B(n1003), .C(n1011), .A(n455), .Y(N13113) );
  OAI21X1 U1472 ( .B(n1004), .C(n1011), .A(n455), .Y(N13104) );
  OAI21X1 U1473 ( .B(n1005), .C(n1011), .A(n455), .Y(N13095) );
  OAI21X1 U1474 ( .B(n1006), .C(n1011), .A(n455), .Y(N13086) );
  OAI21X1 U1475 ( .B(n1000), .C(n1013), .A(n455), .Y(N13077) );
  OAI21X1 U1476 ( .B(n1002), .C(n1013), .A(n455), .Y(N13068) );
  OAI21X1 U1477 ( .B(n2073), .C(n1013), .A(n455), .Y(N13059) );
  OAI21X1 U1478 ( .B(n1661), .C(n1013), .A(n455), .Y(N13050) );
  OAI21X1 U1479 ( .B(n1003), .C(n1013), .A(n455), .Y(N13041) );
  OAI21X1 U1480 ( .B(n1004), .C(n1013), .A(n455), .Y(N13032) );
  OAI21X1 U1481 ( .B(n1005), .C(n1013), .A(n456), .Y(N13023) );
  OAI21X1 U1482 ( .B(n1006), .C(n1013), .A(n456), .Y(N13014) );
  OAI31XL U1483 ( .A(n1245), .B(n440), .C(n438), .D(n463), .Y(N12686) );
  OAI31XL U1484 ( .A(n1245), .B(dps[0]), .C(n440), .D(n463), .Y(N12679) );
  OAI31XL U1485 ( .A(n1245), .B(dps[1]), .C(n438), .D(n463), .Y(N12672) );
  OAI31XL U1486 ( .A(n1247), .B(n440), .C(n438), .D(n463), .Y(N12658) );
  OAI31XL U1487 ( .A(n1247), .B(dps[0]), .C(n440), .D(n463), .Y(N12651) );
  OAI31XL U1488 ( .A(n1247), .B(dps[1]), .C(n438), .D(n463), .Y(N12644) );
  NAND2X1 U1489 ( .A(n1246), .B(n441), .Y(n1247) );
  ENOX1 U1490 ( .A(n117), .B(n1242), .C(dpc[5]), .D(n1243), .Y(N12695) );
  ENOX1 U1491 ( .A(n437), .B(n1242), .C(dpc[3]), .D(n1243), .Y(N12693) );
  ENOX1 U1492 ( .A(n435), .B(n1242), .C(dpc[4]), .D(n1243), .Y(N12694) );
  OAI211X1 U1493 ( .C(n2112), .D(n1808), .A(n463), .B(n486), .Y(N13366) );
  INVX1 U1494 ( .A(n482), .Y(n1939) );
  NAND21X1 U1495 ( .B(n1941), .A(n387), .Y(n482) );
  NAND31X1 U1496 ( .C(n398), .A(n2113), .B(n1735), .Y(n998) );
  NAND32X1 U1497 ( .B(n1840), .C(n398), .A(n1804), .Y(n723) );
  NOR21XL U1498 ( .B(multemp2[2]), .A(n998), .Y(N13325) );
  NOR21XL U1499 ( .B(multemp2[3]), .A(n998), .Y(N13326) );
  NOR21XL U1500 ( .B(multemp2[4]), .A(n998), .Y(N13327) );
  NOR21XL U1501 ( .B(multemp2[5]), .A(n998), .Y(N13328) );
  NOR21XL U1502 ( .B(multemp2[6]), .A(n998), .Y(N13329) );
  NOR21XL U1503 ( .B(multemp2[7]), .A(n998), .Y(N13330) );
  NOR21XL U1504 ( .B(multemp2[8]), .A(n998), .Y(N13331) );
  NOR21XL U1505 ( .B(multemp2[9]), .A(n998), .Y(N13332) );
  NOR21XL U1506 ( .B(n394), .A(n1807), .Y(N10562) );
  NOR4XL U1507 ( .A(n1815), .B(n1816), .C(n1071), .D(n1066), .Y(n1807) );
  OAI211X1 U1508 ( .C(n1940), .D(n1818), .A(n1819), .B(n1820), .Y(n1815) );
  AOI32X1 U1509 ( .A(n1940), .B(n124), .C(n1817), .D(n1765), .E(n1764), .Y(
        n1816) );
  INVX1 U1510 ( .A(pc_i[4]), .Y(n859) );
  INVX1 U1511 ( .A(pc_i[6]), .Y(n941) );
  INVX1 U1512 ( .A(pc_i[5]), .Y(n2061) );
  OR2X1 U1513 ( .A(n458), .B(n173), .Y(N13324) );
  AOI21X1 U1514 ( .B(n2113), .C(n487), .A(n396), .Y(n173) );
  NAND2X1 U1515 ( .A(n1015), .B(n1942), .Y(n1309) );
  AND3X1 U1516 ( .A(n389), .B(n1941), .C(n1460), .Y(N584) );
  AND3X1 U1517 ( .A(n730), .B(n393), .C(n1941), .Y(N585) );
  AND3X1 U1518 ( .A(n389), .B(n1940), .C(n1763), .Y(N12912) );
  AND2X1 U1519 ( .A(sfroe_comb_s), .B(n392), .Y(N11488) );
  INVX1 U1520 ( .A(n955), .Y(sfroe_comb_s) );
  NAND21X1 U1521 ( .B(n1298), .A(n954), .Y(n955) );
  AND2X1 U1522 ( .A(n391), .B(n1299), .Y(N11486) );
  AND2X1 U1523 ( .A(n500), .B(n502), .Y(N13367) );
  INVX1 U1524 ( .A(n1078), .Y(n1840) );
  OAI21X1 U1525 ( .B(n1126), .C(n397), .A(n456), .Y(N12722) );
  NOR4XL U1526 ( .A(n1127), .B(n1128), .C(n22), .D(n2040), .Y(n1126) );
  NAND2X1 U1527 ( .A(n1129), .B(n1109), .Y(n1127) );
  AOI31X1 U1528 ( .A(n1800), .B(n972), .C(n2081), .D(n399), .Y(N10569) );
  NOR2X1 U1529 ( .A(n125), .B(n723), .Y(N680) );
  NOR2X1 U1530 ( .A(n1954), .B(n723), .Y(N683) );
  NOR2X1 U1531 ( .A(n2078), .B(n723), .Y(N682) );
  OR2X1 U1532 ( .A(n459), .B(n174), .Y(n1024) );
  AOI21X1 U1533 ( .B(n7), .C(n1710), .A(n1690), .Y(n174) );
  INVX1 U1534 ( .A(pc_i[2]), .Y(n928) );
  INVX1 U1535 ( .A(pc_i[3]), .Y(n869) );
  AOI21BBXL U1536 ( .B(cpu_resume), .C(irq), .A(n458), .Y(N13379) );
  INVX1 U1537 ( .A(pc_i[7]), .Y(n824) );
  NAND43X1 U1538 ( .B(n475), .C(n474), .D(n459), .A(n473), .Y(N12977) );
  INVX1 U1539 ( .A(n472), .Y(n473) );
  AND3X1 U1540 ( .A(mempsack), .B(n471), .C(n470), .Y(n474) );
  INVX1 U1541 ( .A(n1710), .Y(n475) );
  INVX1 U1542 ( .A(pc_i[0]), .Y(n1197) );
  NOR2X1 U1543 ( .A(n120), .B(n658), .Y(retiinstr) );
  NOR21XL U1544 ( .B(n1351), .A(n1350), .Y(n1568) );
  NAND21X1 U1545 ( .B(n125), .A(n1344), .Y(n1351) );
  AOI21BBXL U1546 ( .B(n977), .C(n978), .A(n429), .Y(n1350) );
  MUX2X1 U1547 ( .D0(N13352), .D1(n189), .S(N13353), .Y(n1607) );
  AO22X1 U1548 ( .A(memdatai[0]), .B(n1072), .C(ramdatai[0]), .D(n1071), .Y(
        n1102) );
  AOI21X1 U1549 ( .B(n725), .C(n2009), .A(n726), .Y(n696) );
  MUX2X1 U1550 ( .D0(N13350), .D1(n187), .S(N13353), .Y(n493) );
  MUX2X1 U1551 ( .D0(N13348), .D1(n185), .S(N13353), .Y(n494) );
  MUX2X1 U1552 ( .D0(N13346), .D1(divtemp1_0_), .S(N13353), .Y(n495) );
  MUX2X1 U1553 ( .D0(N13351), .D1(n188), .S(N13353), .Y(n496) );
  MUX2X1 U1554 ( .D0(N13349), .D1(n186), .S(N13353), .Y(n497) );
  MUX2X1 U1555 ( .D0(N13347), .D1(n184), .S(N13353), .Y(n498) );
  NAND21X1 U1556 ( .B(n1078), .A(n696), .Y(n695) );
  INVX1 U1557 ( .A(n1632), .Y(n775) );
  INVX1 U1558 ( .A(n795), .Y(n1610) );
  INVX1 U1559 ( .A(n1616), .Y(n801) );
  INVX1 U1560 ( .A(n1617), .Y(n790) );
  INVX1 U1561 ( .A(n1621), .Y(n785) );
  INVX1 U1562 ( .A(n1623), .Y(n780) );
  INVX1 U1563 ( .A(pc_i[13]), .Y(n2056) );
  INVX1 U1564 ( .A(n1613), .Y(n812) );
  INVX1 U1565 ( .A(n1615), .Y(n807) );
  INVX1 U1566 ( .A(n1612), .Y(n817) );
  INVX1 U1567 ( .A(n868), .Y(n1903) );
  AND2X1 U1568 ( .A(n1482), .B(n1468), .Y(n1398) );
  INVX1 U1569 ( .A(n1540), .Y(n1482) );
  MUX2X1 U1570 ( .D0(n1966), .D1(n2161), .S(n1571), .Y(n1603) );
  INVX1 U1571 ( .A(n1656), .Y(n842) );
  INVX1 U1572 ( .A(n1655), .Y(n848) );
  INVX1 U1573 ( .A(n1659), .Y(n836) );
  AOI22AXL U1574 ( .A(n1961), .B(n1916), .D(n1470), .C(n1468), .Y(n1384) );
  MUX2IX1 U1575 ( .D0(n2154), .D1(n2152), .S(n1571), .Y(n175) );
  MUX2IX1 U1576 ( .D0(n2140), .D1(n2155), .S(n1571), .Y(n176) );
  INVX1 U1577 ( .A(n1361), .Y(n1912) );
  INVX1 U1578 ( .A(n969), .Y(n1900) );
  INVX1 U1579 ( .A(n726), .Y(n2008) );
  MUX2X1 U1580 ( .D0(n1556), .D1(n1965), .S(n1571), .Y(n1557) );
  INVX1 U1581 ( .A(n1645), .Y(n860) );
  INVX1 U1582 ( .A(n1646), .Y(n854) );
  INVX1 U1583 ( .A(n1644), .Y(n866) );
  MUX2IX1 U1584 ( .D0(n2159), .D1(n2157), .S(n1571), .Y(n177) );
  INVX1 U1585 ( .A(n968), .Y(n1901) );
  INVX1 U1586 ( .A(n967), .Y(n1902) );
  OAI22X1 U1587 ( .A(n1499), .B(n45), .C(n1950), .D(n29), .Y(n1498) );
  NOR4XL U1588 ( .A(multemp2[9]), .B(multemp2[8]), .C(multemp2[7]), .D(
        multemp2[6]), .Y(n1175) );
  MUX2X1 U1589 ( .D0(n1967), .D1(n1964), .S(n1571), .Y(n1330) );
  INVX1 U1590 ( .A(n1642), .Y(n926) );
  INVX1 U1591 ( .A(n1643), .Y(n872) );
  NOR21XL U1592 ( .B(n658), .A(n1136), .Y(n1129) );
  INVX1 U1593 ( .A(pc_i[15]), .Y(n2054) );
  INVX1 U1594 ( .A(pc_i[14]), .Y(n2055) );
  INVX1 U1595 ( .A(n1323), .Y(n1981) );
  OAI221X1 U1596 ( .A(n2060), .B(n77), .C(n1267), .D(n31), .E(n1324), .Y(n1323) );
  INVX1 U1597 ( .A(pc_i[8]), .Y(n2060) );
  AOI222XL U1598 ( .A(N11786), .B(n1269), .C(N11820), .D(n1270), .E(N11803), 
        .F(n1271), .Y(n1324) );
  INVX1 U1599 ( .A(n1286), .Y(n1988) );
  OAI221X1 U1600 ( .A(n987), .B(n77), .C(n1267), .D(n43), .E(n1287), .Y(n1286)
         );
  AOI222XL U1601 ( .A(n43), .B(n1269), .C(n43), .D(n98), .E(N11796), .F(n111), 
        .Y(n1287) );
  INVX1 U1602 ( .A(n1284), .Y(n1987) );
  OAI221X1 U1603 ( .A(n928), .B(n77), .C(n1267), .D(n33), .E(n1285), .Y(n1284)
         );
  AOI222XL U1604 ( .A(N11780), .B(n1269), .C(N11814), .D(n1270), .E(N11797), 
        .F(n1271), .Y(n1285) );
  INVX1 U1605 ( .A(n1282), .Y(n1986) );
  OAI221X1 U1606 ( .A(n869), .B(n77), .C(n1267), .D(n45), .E(n1283), .Y(n1282)
         );
  AOI222XL U1607 ( .A(N11781), .B(n1269), .C(N11815), .D(n98), .E(N11798), .F(
        n111), .Y(n1283) );
  INVX1 U1608 ( .A(n1280), .Y(n1985) );
  OAI221X1 U1609 ( .A(n859), .B(n77), .C(n1267), .D(n53), .E(n1281), .Y(n1280)
         );
  AOI222XL U1610 ( .A(N11782), .B(n1269), .C(N11816), .D(n1270), .E(N11799), 
        .F(n1271), .Y(n1281) );
  INVX1 U1611 ( .A(n1276), .Y(n1983) );
  OAI221X1 U1612 ( .A(n941), .B(n77), .C(n1267), .D(n25), .E(n1277), .Y(n1276)
         );
  AOI222XL U1613 ( .A(N11784), .B(n1269), .C(N11818), .D(n98), .E(N11801), .F(
        n111), .Y(n1277) );
  INVX1 U1614 ( .A(n1265), .Y(n1982) );
  OAI221X1 U1615 ( .A(n824), .B(n77), .C(n1267), .D(n50), .E(n1268), .Y(n1265)
         );
  AOI222XL U1616 ( .A(N11785), .B(n1269), .C(N11819), .D(n1270), .E(N11802), 
        .F(n1271), .Y(n1268) );
  INVX1 U1617 ( .A(n1320), .Y(n1980) );
  OAI221X1 U1618 ( .A(n984), .B(n77), .C(n1267), .D(n39), .E(n1321), .Y(n1320)
         );
  AOI222XL U1619 ( .A(N11787), .B(n1269), .C(N11821), .D(n98), .E(N11804), .F(
        n111), .Y(n1321) );
  NOR4XL U1620 ( .A(multemp2[5]), .B(multemp2[4]), .C(multemp2[3]), .D(
        multemp2[2]), .Y(n1174) );
  INVX1 U1621 ( .A(n1132), .Y(n2022) );
  NOR32XL U1622 ( .B(n1105), .C(n1069), .A(n1106), .Y(n1089) );
  NOR32XL U1623 ( .B(n1194), .C(n1195), .A(n1178), .Y(n1187) );
  INVX1 U1624 ( .A(N11555), .Y(n2063) );
  INVX1 U1625 ( .A(pc_i[11]), .Y(n2058) );
  INVX1 U1626 ( .A(pc_i[12]), .Y(n2057) );
  AND3X1 U1627 ( .A(n1103), .B(n1104), .C(n2090), .Y(n1108) );
  AND2X1 U1628 ( .A(n1108), .B(n1109), .Y(n1105) );
  NAND3X1 U1629 ( .A(n1129), .B(n1109), .C(n1128), .Y(n1138) );
  NAND3X1 U1630 ( .A(n2025), .B(n1151), .C(n1129), .Y(n1134) );
  INVX1 U1631 ( .A(dpc[1]), .Y(n2164) );
  INVX1 U1632 ( .A(dpc[2]), .Y(n2165) );
  NAND3X1 U1633 ( .A(dpc[1]), .B(dpc[0]), .C(dpc[2]), .Y(n1326) );
  INVX1 U1634 ( .A(n1136), .Y(n2021) );
  NAND3X1 U1635 ( .A(dpc[0]), .B(n2165), .C(dpc[1]), .Y(n1325) );
  NAND3X1 U1636 ( .A(dpc[0]), .B(n2164), .C(dpc[2]), .Y(n1327) );
  NAND3X1 U1637 ( .A(n2164), .B(n2165), .C(dpc[0]), .Y(n1329) );
  NAND4X1 U1638 ( .A(n1123), .B(n446), .C(n69), .D(n89), .Y(n1122) );
  NOR21XL U1639 ( .B(n1103), .A(n1104), .Y(n1070) );
  AND4X1 U1640 ( .A(n1356), .B(n1196), .C(n1226), .D(n92), .Y(n1195) );
  NOR2X1 U1641 ( .A(n2091), .B(n124), .Y(n1066) );
  INVX1 U1642 ( .A(pc_i[10]), .Y(n2059) );
  INVX1 U1643 ( .A(n1183), .Y(n1925) );
  AND3X1 U1644 ( .A(n118), .B(n437), .C(n434), .Y(n178) );
  OAI22X1 U1645 ( .A(n33), .B(n1094), .C(n2059), .D(n1069), .Y(n1093) );
  NAND4X1 U1646 ( .A(n1194), .B(n1951), .C(n1195), .D(n1355), .Y(n1348) );
  AOI221XL U1647 ( .A(n1926), .B(n2113), .C(n1925), .D(n2112), .E(n2046), .Y(
        n1355) );
  NOR3XL U1648 ( .A(n2102), .B(n57), .C(n2033), .Y(n1766) );
  INVX1 U1649 ( .A(n991), .Y(n1889) );
  NAND32X1 U1650 ( .B(n1821), .C(n56), .A(n912), .Y(n991) );
  INVX1 U1651 ( .A(n1109), .Y(n2025) );
  AND3X1 U1652 ( .A(n119), .B(n435), .C(n436), .Y(n179) );
  AND3X1 U1653 ( .A(n434), .B(n119), .C(n436), .Y(n180) );
  AND3X1 U1654 ( .A(n435), .B(n437), .C(n118), .Y(n181) );
  OR2X1 U1655 ( .A(n885), .B(n2078), .Y(n1107) );
  INVX1 U1656 ( .A(n1151), .Y(n2040) );
  NAND43X1 U1657 ( .B(n16), .C(n445), .D(n2100), .A(n1597), .Y(n1803) );
  AND2X1 U1658 ( .A(n1740), .B(n1922), .Y(n1797) );
  AND3X1 U1659 ( .A(n733), .B(n734), .C(n1945), .Y(n730) );
  OAI21X1 U1660 ( .B(n120), .C(n56), .A(n737), .Y(n733) );
  OAI22X1 U1661 ( .A(n2068), .B(n2077), .C(n125), .D(n736), .Y(n734) );
  NOR2X1 U1662 ( .A(n2096), .B(n2089), .Y(n1792) );
  NAND2X1 U1663 ( .A(n1609), .B(n1839), .Y(n1779) );
  NAND2X1 U1664 ( .A(n1598), .B(n1118), .Y(n1775) );
  NAND2X1 U1665 ( .A(n1822), .B(n1946), .Y(n1800) );
  INVX1 U1666 ( .A(n1347), .Y(n1949) );
  NAND2X1 U1667 ( .A(n1740), .B(n902), .Y(n1770) );
  NAND2X1 U1668 ( .A(n1598), .B(n1686), .Y(n1774) );
  NAND2X1 U1669 ( .A(n1737), .B(n902), .Y(n1769) );
  NAND2X1 U1670 ( .A(n1910), .B(n1839), .Y(n1780) );
  OR2X1 U1671 ( .A(n897), .B(n449), .Y(n1765) );
  INVX1 U1672 ( .A(n1069), .Y(n1095) );
  OAI22X1 U1673 ( .A(n2141), .B(n1030), .C(n2142), .D(n1029), .Y(N12970) );
  OAI22X1 U1674 ( .A(n2136), .B(n1030), .C(n2138), .D(n1029), .Y(N12971) );
  OAI22X1 U1675 ( .A(n2134), .B(n1030), .C(n2135), .D(n1029), .Y(N12969) );
  OAI22X1 U1676 ( .A(n2053), .B(n1030), .C(n2125), .D(n1029), .Y(N12965) );
  OAI22X1 U1677 ( .A(n2064), .B(n1030), .C(n2124), .D(n1029), .Y(N12966) );
  OAI22X1 U1678 ( .A(n2120), .B(n1030), .C(n2123), .D(n1029), .Y(N12967) );
  NOR2X1 U1679 ( .A(rst), .B(n1031), .Y(N12968) );
  INVX1 U1680 ( .A(n1014), .Y(n2073) );
  INVX1 U1681 ( .A(n680), .Y(n1291) );
  NAND21X1 U1682 ( .B(n1941), .A(n730), .Y(n1469) );
  INVX1 U1683 ( .A(n684), .Y(cs_run) );
  INVX1 U1684 ( .A(n1562), .Y(n677) );
  AO21X1 U1685 ( .B(n1424), .C(pc_o[9]), .A(n740), .Y(n762) );
  OAI22X1 U1686 ( .A(n1458), .B(n984), .C(n1457), .D(n987), .Y(n761) );
  OAI21AX1 U1687 ( .B(sfroe_r), .C(sfrwe_r), .A(sfrack), .Y(n471) );
  AND3X2 U1688 ( .A(n738), .B(n1953), .C(n182), .Y(n1292) );
  NOR32XL U1689 ( .B(n653), .C(n112), .A(n1131), .Y(n698) );
  NAND21X1 U1690 ( .B(n665), .A(n664), .Y(n697) );
  MUX2X1 U1691 ( .D0(n219), .D1(n218), .S(n244), .Y(dph[6]) );
  MUX4X1 U1692 ( .D0(dph_reg[6]), .D1(dph_reg[14]), .D2(dph_reg[22]), .D3(
        dph_reg[30]), .S0(n250), .S1(n246), .Y(n219) );
  MUX4X1 U1693 ( .D0(dph_reg[38]), .D1(dph_reg[46]), .D2(dph_reg[54]), .D3(
        dph_reg[62]), .S0(n250), .S1(n246), .Y(n218) );
  NOR21XL U1694 ( .B(c), .A(n666), .Y(n692) );
  MUX2X1 U1695 ( .D0(n217), .D1(n216), .S(n244), .Y(dph[7]) );
  MUX2X1 U1696 ( .D0(n201), .D1(n200), .S(dps[2]), .Y(dpl[7]) );
  MUX2X1 U1697 ( .D0(n203), .D1(n202), .S(dps[2]), .Y(dpl[6]) );
  MUX4X1 U1698 ( .D0(dpl_reg[6]), .D1(dpl_reg[14]), .D2(dpl_reg[22]), .D3(
        dpl_reg[30]), .S0(n249), .S1(dps[1]), .Y(n203) );
  MUX2X1 U1699 ( .D0(n231), .D1(n230), .S(n245), .Y(dph[0]) );
  MUX4X1 U1700 ( .D0(dph_reg[0]), .D1(dph_reg[8]), .D2(dph_reg[16]), .D3(
        dph_reg[24]), .S0(n251), .S1(n247), .Y(n231) );
  MUX4X1 U1701 ( .D0(dph_reg[32]), .D1(dph_reg[40]), .D2(dph_reg[48]), .D3(
        dph_reg[56]), .S0(n251), .S1(n247), .Y(n230) );
  MUX2X1 U1702 ( .D0(n221), .D1(n220), .S(n244), .Y(dph[5]) );
  MUX4X1 U1703 ( .D0(dph_reg[5]), .D1(dph_reg[13]), .D2(dph_reg[21]), .D3(
        dph_reg[29]), .S0(n250), .S1(n246), .Y(n221) );
  MUX4X1 U1704 ( .D0(dph_reg[37]), .D1(dph_reg[45]), .D2(dph_reg[53]), .D3(
        dph_reg[61]), .S0(n250), .S1(n246), .Y(n220) );
  MUX2X1 U1705 ( .D0(n223), .D1(n222), .S(n244), .Y(dph[4]) );
  MUX4X1 U1706 ( .D0(dph_reg[4]), .D1(dph_reg[12]), .D2(dph_reg[20]), .D3(
        dph_reg[28]), .S0(n250), .S1(n246), .Y(n223) );
  MUX4X1 U1707 ( .D0(dph_reg[36]), .D1(dph_reg[44]), .D2(dph_reg[52]), .D3(
        dph_reg[60]), .S0(n250), .S1(n246), .Y(n222) );
  MUX2X1 U1708 ( .D0(n209), .D1(n208), .S(n244), .Y(dpl[3]) );
  MUX4X1 U1709 ( .D0(dpl_reg[3]), .D1(dpl_reg[11]), .D2(dpl_reg[19]), .D3(
        dpl_reg[27]), .S0(dps[0]), .S1(N350), .Y(n209) );
  MUX2X1 U1710 ( .D0(n213), .D1(n212), .S(n244), .Y(dpl[1]) );
  MUX4X1 U1711 ( .D0(dpl_reg[1]), .D1(dpl_reg[9]), .D2(dpl_reg[17]), .D3(
        dpl_reg[25]), .S0(n249), .S1(N350), .Y(n213) );
  MUX2X1 U1712 ( .D0(n215), .D1(n214), .S(n244), .Y(dpl[0]) );
  MUX4X1 U1713 ( .D0(dpl_reg[0]), .D1(dpl_reg[8]), .D2(dpl_reg[16]), .D3(
        dpl_reg[24]), .S0(n250), .S1(n246), .Y(n215) );
  MUX4X1 U1714 ( .D0(dpl_reg[32]), .D1(dpl_reg[40]), .D2(dpl_reg[48]), .D3(
        dpl_reg[56]), .S0(n250), .S1(n246), .Y(n214) );
  MUX2X1 U1715 ( .D0(n205), .D1(n204), .S(n244), .Y(dpl[5]) );
  MUX4X1 U1716 ( .D0(dpl_reg[5]), .D1(dpl_reg[13]), .D2(dpl_reg[21]), .D3(
        dpl_reg[29]), .S0(n249), .S1(N350), .Y(n205) );
  MUX4X1 U1717 ( .D0(dpl_reg[37]), .D1(dpl_reg[45]), .D2(dpl_reg[53]), .D3(
        dpl_reg[61]), .S0(n249), .S1(N350), .Y(n204) );
  MUX2X1 U1718 ( .D0(n207), .D1(n206), .S(n244), .Y(dpl[4]) );
  MUX4X1 U1719 ( .D0(dpl_reg[4]), .D1(dpl_reg[12]), .D2(dpl_reg[20]), .D3(
        dpl_reg[28]), .S0(n249), .S1(dps[1]), .Y(n207) );
  MUX4X1 U1720 ( .D0(dpl_reg[36]), .D1(dpl_reg[44]), .D2(dpl_reg[52]), .D3(
        dpl_reg[60]), .S0(n249), .S1(N350), .Y(n206) );
  AO2222XL U1721 ( .A(n957), .B(pc_i[11]), .C(n956), .D(temp[3]), .E(
        alu_out[11]), .F(n1160), .G(n384), .H(n1616), .Y(n876) );
  MUX2X1 U1722 ( .D0(pc_o[11]), .D1(n1502), .S(n451), .Y(memaddr_comb[11]) );
  MUX2BXL U1723 ( .D0(memrd), .D1(n1461), .S(n450), .Y(memrd_comb) );
  NAND21X1 U1724 ( .B(n2072), .A(n1460), .Y(n1461) );
  MUX2X1 U1725 ( .D0(n49), .D1(n1504), .S(n450), .Y(memaddr_comb[13]) );
  AO2222XL U1726 ( .A(n957), .B(pc_i[12]), .C(n956), .D(temp[4]), .E(
        alu_out[12]), .F(n113), .G(n384), .H(n1617), .Y(n867) );
  AO2222XL U1727 ( .A(n957), .B(pc_i[13]), .C(n956), .D(temp[5]), .E(
        alu_out[13]), .F(n1160), .G(n384), .H(n1621), .Y(n858) );
  AO2222XL U1728 ( .A(n957), .B(pc_i[14]), .C(n956), .D(temp[6]), .E(
        alu_out[14]), .F(n113), .G(n384), .H(n1623), .Y(n850) );
  MUX2X1 U1729 ( .D0(pc_o[14]), .D1(n1505), .S(waitstaten), .Y(
        memaddr_comb[14]) );
  MUX2X1 U1730 ( .D0(pc_o[12]), .D1(n1503), .S(waitstaten), .Y(
        memaddr_comb[12]) );
  MUX2BXL U1731 ( .D0(ramwe), .D1(n183), .S(n451), .Y(ramwe_comb) );
  AOI21X1 U1732 ( .B(n1298), .C(n1297), .A(n1296), .Y(n183) );
  MUX2X1 U1733 ( .D0(ramoe), .D1(n1299), .S(n450), .Y(ramoe_comb) );
  MUX2X1 U1734 ( .D0(mempsrd), .D1(n1474), .S(waitstaten), .Y(mempsrd_comb) );
  AO2222XL U1735 ( .A(n957), .B(pc_i[15]), .C(n956), .D(temp[7]), .E(
        alu_out[15]), .F(n1160), .G(n384), .H(n1632), .Y(n961) );
  MUX2X1 U1736 ( .D0(pc_o[15]), .D1(n1632), .S(n86), .Y(N12856) );
  MUX2X1 U1737 ( .D0(n1361), .D1(temp[2]), .S(n808), .Y(N12826) );
  MUX2X1 U1738 ( .D0(memaddr[2]), .D1(n1644), .S(n622), .Y(N12843) );
  MUX2X1 U1739 ( .D0(n868), .D1(temp[3]), .S(n808), .Y(N12827) );
  MUX2X1 U1740 ( .D0(memaddr[3]), .D1(n1645), .S(n622), .Y(N12844) );
  MUX2X1 U1741 ( .D0(n967), .D1(temp[4]), .S(n808), .Y(N12828) );
  MUX2X1 U1742 ( .D0(memaddr[4]), .D1(n1646), .S(n622), .Y(N12845) );
  MUX2X1 U1743 ( .D0(n968), .D1(temp[5]), .S(n808), .Y(N12829) );
  MUX2X1 U1744 ( .D0(memaddr[5]), .D1(n1655), .S(n622), .Y(N12846) );
  MUX2X1 U1745 ( .D0(n964), .D1(temp[1]), .S(n808), .Y(N12825) );
  MUX2X1 U1746 ( .D0(memaddr[1]), .D1(n1643), .S(n622), .Y(N12842) );
  NAND43X1 U1747 ( .B(n551), .C(n550), .D(n549), .A(n548), .Y(n963) );
  OAI22X1 U1748 ( .A(n560), .B(n2140), .C(n2133), .D(n541), .Y(n551) );
  OAI221X1 U1749 ( .A(n2127), .B(n2048), .C(n545), .D(n544), .E(n543), .Y(n550) );
  AO21X1 U1750 ( .B(n1926), .C(acc[2]), .A(n547), .Y(n549) );
  OAI31XL U1751 ( .A(n803), .B(n802), .C(n800), .D(n799), .Y(n806) );
  MUX2X1 U1752 ( .D0(n792), .D1(n910), .S(n789), .Y(n800) );
  AO222X1 U1753 ( .A(n1759), .B(phase[2]), .C(n798), .D(n432), .E(n1027), .F(
        phase[3]), .Y(n799) );
  AOI31X1 U1754 ( .A(n794), .B(n781), .C(n885), .D(n779), .Y(n802) );
  MUX2X1 U1755 ( .D0(pc_o[15]), .D1(n1506), .S(n451), .Y(memaddr_comb[15]) );
  MUX2X1 U1756 ( .D0(n969), .D1(temp[6]), .S(n808), .Y(N12830) );
  MUX2X1 U1757 ( .D0(pc_o[6]), .D1(n1656), .S(n622), .Y(N12847) );
  MUX2X1 U1758 ( .D0(n963), .D1(temp[0]), .S(n808), .Y(N12824) );
  NAND21X1 U1759 ( .B(n935), .A(n934), .Y(n1478) );
  AO2222XL U1760 ( .A(alu_out[2]), .B(n113), .C(n385), .D(n1644), .E(n1897), 
        .F(n2015), .G(n1896), .H(ramdatai[2]), .Y(n935) );
  OA2222XL U1761 ( .A(n1202), .B(n2162), .C(n1993), .D(n1198), .E(n928), .F(
        n1193), .G(n33), .H(n1161), .Y(n934) );
  NAND21X1 U1762 ( .B(n862), .A(n861), .Y(n1481) );
  AO2222XL U1763 ( .A(alu_out[4]), .B(n1160), .C(n385), .D(n1646), .E(n1897), 
        .F(n2013), .G(n1896), .H(ramdatai[4]), .Y(n862) );
  OA2222XL U1764 ( .A(n1202), .B(n2156), .C(n1996), .D(n1198), .E(n1193), .F(
        n859), .G(n53), .H(n1161), .Y(n861) );
  NAND21X1 U1765 ( .B(n943), .A(n942), .Y(n1484) );
  OA2222XL U1766 ( .A(n1202), .B(n2139), .C(n1998), .D(n1198), .E(n1193), .F(
        n941), .G(n25), .H(n1161), .Y(n942) );
  AO2222XL U1767 ( .A(alu_out[6]), .B(n113), .C(n385), .D(n1656), .E(n1897), 
        .F(n2011), .G(n1896), .H(ramdatai[6]), .Y(n943) );
  NAND21X1 U1768 ( .B(n855), .A(n852), .Y(n1483) );
  OA2222XL U1769 ( .A(n1202), .B(n2158), .C(n1997), .D(n1198), .E(n2061), .F(
        n1193), .G(n23), .H(n1161), .Y(n852) );
  AO2222XL U1770 ( .A(alu_out[5]), .B(n1160), .C(n385), .D(n1655), .E(n1897), 
        .F(n2012), .G(n1896), .H(ramdatai[5]), .Y(n855) );
  OAI211X1 U1771 ( .C(n948), .D(n1455), .A(n947), .B(n658), .Y(n1299) );
  NAND32X1 U1772 ( .B(n125), .C(instr[3]), .A(n1691), .Y(n947) );
  INVX1 U1773 ( .A(n954), .Y(n948) );
  OAI211X1 U1774 ( .C(n1692), .D(n69), .A(n1693), .B(n1694), .Y(n1691) );
  INVX1 U1775 ( .A(n485), .Y(divtemp1_0_) );
  MUX2AXL U1776 ( .D0(N13336), .D1(n1966), .S(N13343), .Y(n485) );
  MUX2X1 U1777 ( .D0(N13337), .D1(divtempreg[0]), .S(N13343), .Y(n184) );
  MUX2X1 U1778 ( .D0(pc_o[8]), .D1(n1612), .S(n622), .Y(N12849) );
  MUX2X1 U1779 ( .D0(memaddr[9]), .D1(n1613), .S(n622), .Y(N12850) );
  MUX2X1 U1780 ( .D0(pc_o[7]), .D1(n1659), .S(n622), .Y(N12848) );
  AO21X1 U1781 ( .B(n603), .C(n970), .A(n1894), .Y(N12831) );
  MUX2X1 U1782 ( .D0(pc_o[10]), .D1(n1615), .S(n86), .Y(N12851) );
  MUX2X1 U1783 ( .D0(pc_o[11]), .D1(n1616), .S(n86), .Y(N12852) );
  MUX2X1 U1784 ( .D0(pc_o[12]), .D1(n1617), .S(n86), .Y(N12853) );
  MUX2X1 U1785 ( .D0(n49), .D1(n1621), .S(n86), .Y(N12854) );
  MUX2X1 U1786 ( .D0(pc_o[14]), .D1(n1623), .S(n86), .Y(N12855) );
  NAND21X1 U1787 ( .B(n873), .A(n870), .Y(n1479) );
  AO2222XL U1788 ( .A(alu_out[3]), .B(n113), .C(n385), .D(n1645), .E(n1896), 
        .F(ramdatai[3]), .G(n1897), .H(n2014), .Y(n873) );
  OA2222XL U1789 ( .A(n1202), .B(n2153), .C(n1995), .D(n1198), .E(n1193), .F(
        n869), .G(n45), .H(n1161), .Y(n870) );
  NAND21X1 U1790 ( .B(n826), .A(n825), .Y(n1485) );
  OA2222XL U1791 ( .A(n1202), .B(n2160), .C(n1999), .D(n1198), .E(n1193), .F(
        n824), .G(n50), .H(n1161), .Y(n825) );
  AO2222XL U1792 ( .A(alu_out[7]), .B(n1160), .C(n385), .D(n1659), .E(n1896), 
        .F(ramdatai[7]), .G(n1897), .H(n2010), .Y(n826) );
  NAND21X1 U1793 ( .B(n879), .A(n878), .Y(n1501) );
  OA2222XL U1794 ( .A(n27), .B(n976), .C(n1964), .D(n975), .E(n2120), .F(n974), 
        .G(n2148), .H(n973), .Y(n878) );
  AO2222XL U1795 ( .A(n384), .B(n1615), .C(n971), .D(pc_i[10]), .E(n1898), .F(
        instr[7]), .G(alu_out[10]), .H(n113), .Y(n879) );
  NAND21X1 U1796 ( .B(n927), .A(n925), .Y(n1500) );
  OA2222XL U1797 ( .A(n39), .B(n976), .C(n2151), .D(n975), .E(n2064), .F(n974), 
        .G(n2149), .H(n973), .Y(n925) );
  AO2222XL U1798 ( .A(n384), .B(n1613), .C(n971), .D(pc_i[9]), .E(n1898), .F(
        n2189), .G(alu_out[9]), .H(n1160), .Y(n927) );
  MUX2X1 U1799 ( .D0(N13338), .D1(divtempreg[1]), .S(N13343), .Y(n185) );
  XNOR2XL U1800 ( .A(acc[3]), .B(n1370), .Y(N11544) );
  OAI21X1 U1801 ( .B(n1372), .C(n2153), .A(n1379), .Y(N11525) );
  XNOR2XL U1802 ( .A(acc[2]), .B(n1370), .Y(N11543) );
  OAI21X1 U1803 ( .B(n1372), .C(n2162), .A(n2107), .Y(N11524) );
  OAI221X1 U1804 ( .A(n2111), .B(n1381), .C(n1372), .D(n1225), .E(n1379), .Y(
        N11522) );
  AOI21BBXL U1805 ( .B(n1539), .C(n1091), .A(n638), .Y(n705) );
  NOR21XL U1806 ( .B(N1761), .A(n644), .Y(n638) );
  AOI222XL U1807 ( .A(n1199), .B(n1200), .C(n770), .D(acc[7]), .E(acc[0]), .F(
        n769), .Y(n771) );
  XNOR2XL U1808 ( .A(n1184), .B(n1229), .Y(n1199) );
  NAND2X1 U1809 ( .A(n2115), .B(n2116), .Y(n1229) );
  AND4X1 U1810 ( .A(n1427), .B(n1428), .C(n1429), .D(n1430), .Y(n670) );
  AOI22X1 U1811 ( .A(pc_o[14]), .B(n1424), .C(pc_o[6]), .D(n22), .Y(n1427) );
  AOI222XL U1812 ( .A(N1767), .B(n1423), .C(temp2_comb[6]), .D(n1909), .E(
        pc_i[14]), .F(n1905), .Y(n1428) );
  AOI222XL U1813 ( .A(n702), .B(n1431), .C(ramdatai[6]), .D(n2079), .E(n969), 
        .F(n1398), .Y(n1430) );
  AND4X1 U1814 ( .A(n1392), .B(n1393), .C(n1394), .D(n1395), .Y(n667) );
  AOI22X1 U1815 ( .A(pc_o[15]), .B(n1424), .C(pc_o[7]), .D(n21), .Y(n1392) );
  AOI222XL U1816 ( .A(N1768), .B(n1423), .C(temp2_comb[7]), .D(n1909), .E(
        pc_i[15]), .F(n1905), .Y(n1393) );
  AOI222XL U1817 ( .A(n702), .B(n1397), .C(ramdatai[7]), .D(n2079), .E(n1398), 
        .F(n970), .Y(n1395) );
  NAND3X1 U1818 ( .A(dec_accop[6]), .B(n2111), .C(n2114), .Y(n1379) );
  OAI211X1 U1819 ( .C(n1885), .D(n1083), .A(n1082), .B(n1079), .Y(n1474) );
  OAI211X1 U1820 ( .C(n742), .D(n743), .A(cs_run), .B(n102), .Y(n1082) );
  AOI31X1 U1821 ( .A(n2008), .B(n725), .C(n1840), .D(n744), .Y(n1083) );
  MUX2X1 U1822 ( .D0(N13339), .D1(divtempreg[2]), .S(N13343), .Y(n186) );
  MUX2X1 U1823 ( .D0(N13340), .D1(divtempreg[3]), .S(N13343), .Y(n187) );
  NOR2X1 U1824 ( .A(dec_accop[8]), .B(dec_accop[10]), .Y(n1371) );
  NAND42X1 U1825 ( .C(dec_accop[18]), .D(dec_accop[16]), .A(n2111), .B(n1405), 
        .Y(n1370) );
  NOR3XL U1826 ( .A(dec_accop[6]), .B(dec_accop[8]), .C(dec_accop[7]), .Y(
        n1405) );
  AOI21BBXL U1827 ( .B(dec_accop[5]), .C(dec_accop[18]), .A(n1381), .Y(n1372)
         );
  XNOR2XL U1828 ( .A(acc[0]), .B(n1370), .Y(N11541) );
  AOI222XL U1829 ( .A(n1919), .B(acc[3]), .C(n1403), .D(n607), .E(n1917), .F(
        n1966), .Y(n594) );
  XNOR2XL U1830 ( .A(n1231), .B(n1232), .Y(n1403) );
  INVX1 U1831 ( .A(n1380), .Y(n2107) );
  GEN2XL U1832 ( .D(acc[3]), .E(n1378), .C(ac), .B(n2108), .A(n2110), .Y(n1380) );
  INVX1 U1833 ( .A(n1375), .Y(n2108) );
  INVX1 U1834 ( .A(acc[1]), .Y(n2127) );
  INVX1 U1835 ( .A(acc[2]), .Y(n1967) );
  INVX1 U1836 ( .A(c), .Y(n2133) );
  NAND3X1 U1837 ( .A(dec_accop[18]), .B(n2111), .C(n2114), .Y(n1375) );
  MUX2X1 U1838 ( .D0(N13341), .D1(divtempreg[4]), .S(N13343), .Y(n188) );
  INVX1 U1839 ( .A(dec_accop[9]), .Y(n2115) );
  INVX1 U1840 ( .A(dec_accop[5]), .Y(n2111) );
  INVX1 U1841 ( .A(n1441), .Y(n671) );
  NAND41X1 U1842 ( .D(n1440), .A(n1448), .B(n1447), .C(n1439), .Y(n1441) );
  AOI222XL U1843 ( .A(memaddr[5]), .B(n22), .C(N1766), .D(n1423), .E(n49), .F(
        n1424), .Y(n1447) );
  AOI31X1 U1844 ( .A(n1421), .B(n1587), .C(n1420), .D(n1432), .Y(n1440) );
  AO222X1 U1845 ( .A(dpl_current[1]), .B(n621), .C(dptr_inc[1]), .D(n620), .E(
        n619), .F(temp[1]), .Y(n1643) );
  ENOX1 U1846 ( .A(n2053), .B(n1275), .C(N11842), .D(n1275), .Y(dpl_current[0]) );
  MUX2X1 U1847 ( .D0(n270), .D1(n269), .S(N348), .Y(N11842) );
  MUX4X1 U1848 ( .D0(dpl_reg[0]), .D1(dpl_reg[8]), .D2(dpl_reg[16]), .D3(
        dpl_reg[24]), .S0(n285), .S1(n287), .Y(n270) );
  MUX4X1 U1849 ( .D0(dpl_reg[32]), .D1(dpl_reg[40]), .D2(dpl_reg[48]), .D3(
        dpl_reg[56]), .S0(n285), .S1(n287), .Y(n269) );
  NAND32X1 U1850 ( .B(n593), .C(n592), .A(n591), .Y(n969) );
  OA22X1 U1851 ( .A(n2136), .B(n92), .C(n1183), .D(n2140), .Y(n591) );
  AO21X1 U1852 ( .B(multemp1_0_), .C(n1926), .A(n1435), .Y(n593) );
  AO2222XL U1853 ( .A(n1556), .B(n1917), .C(adder_out[6]), .D(n607), .E(acc[5]), .F(n590), .G(n1919), .H(acc[2]), .Y(n592) );
  NAND32X1 U1854 ( .B(ramsfraddr[5]), .C(ramsfraddr[6]), .A(n831), .Y(n1663)
         );
  MUX2X1 U1855 ( .D0(ramdatao[3]), .D1(n1401), .S(n451), .Y(ramdatao_comb[3])
         );
  AOI22X1 U1856 ( .A(n2067), .B(ramdatao[3]), .C(n1168), .D(rs[0]), .Y(n1189)
         );
  XNOR2XL U1857 ( .A(acc[1]), .B(n1370), .Y(N11542) );
  MUX2AXL U1858 ( .D0(n1490), .D1(n1684), .S(n1904), .Y(n1401) );
  AND3X1 U1859 ( .A(n1495), .B(n1496), .C(n1497), .Y(n1490) );
  AOI22X1 U1860 ( .A(pc_i[3]), .B(n1906), .C(temp2_comb[3]), .D(n1909), .Y(
        n1495) );
  AOI221XL U1861 ( .A(pc_i[11]), .B(n1905), .C(N1764), .D(n1423), .E(n1498), 
        .Y(n1497) );
  NOR3XL U1862 ( .A(ramsfraddr[0]), .B(ramsfraddr[2]), .C(n2119), .Y(n1014) );
  INVX1 U1863 ( .A(ramsfraddr[1]), .Y(n2119) );
  INVX1 U1864 ( .A(ramsfraddr[4]), .Y(n2163) );
  INVX1 U1865 ( .A(ramsfraddr[0]), .Y(n2071) );
  INVX1 U1866 ( .A(ramsfraddr[2]), .Y(n2121) );
  NOR2X1 U1867 ( .A(n2163), .B(ramsfraddr[3]), .Y(n1012) );
  ENOX1 U1868 ( .A(n2064), .B(n91), .C(N11841), .D(n91), .Y(dpl_current[1]) );
  MUX2X1 U1869 ( .D0(n272), .D1(n271), .S(n118), .Y(N11841) );
  MUX4X1 U1870 ( .D0(dpl_reg[1]), .D1(dpl_reg[9]), .D2(dpl_reg[17]), .D3(
        dpl_reg[25]), .S0(n285), .S1(n287), .Y(n272) );
  MUX4X1 U1871 ( .D0(dpl_reg[33]), .D1(dpl_reg[41]), .D2(dpl_reg[49]), .D3(
        dpl_reg[57]), .S0(n285), .S1(n287), .Y(n271) );
  INVX1 U1872 ( .A(ramsfraddr[7]), .Y(n1961) );
  INVX1 U1873 ( .A(n477), .Y(n831) );
  NAND21X1 U1874 ( .B(n1961), .A(ramsfrwe), .Y(n477) );
  MUX2X1 U1875 ( .D0(N13342), .D1(divtempreg[5]), .S(N13343), .Y(n189) );
  OAI221X1 U1876 ( .A(n1335), .B(n440), .C(n1189), .D(n1336), .E(n1337), .Y(
        N347) );
  AOI32X1 U1877 ( .A(n2074), .B(n2075), .C(ramdatao[1]), .D(n1338), .E(rs[0]), 
        .Y(n1337) );
  OR2X1 U1878 ( .A(dps[3]), .B(n2074), .Y(n1335) );
  INVX1 U1879 ( .A(n1417), .Y(n672) );
  NAND41X1 U1880 ( .D(n1416), .A(n1473), .B(n1471), .C(n1472), .Y(n1417) );
  AOI222XL U1881 ( .A(pc_o[4]), .B(n21), .C(N1765), .D(n1423), .E(pc_o[12]), 
        .F(n1424), .Y(n1473) );
  AOI222XL U1882 ( .A(pc_i[12]), .B(n1905), .C(pc_i[4]), .D(n1906), .E(
        temp2_comb[4]), .F(n1909), .Y(n1471) );
  AO222X1 U1883 ( .A(n619), .B(temp[3]), .C(dptr_inc[3]), .D(n620), .E(n621), 
        .F(dpl_current[3]), .Y(n1645) );
  AO222X1 U1884 ( .A(n619), .B(temp[4]), .C(dptr_inc[4]), .D(n620), .E(n621), 
        .F(dpl_current[4]), .Y(n1646) );
  AO222X1 U1885 ( .A(dpl_current[2]), .B(n621), .C(dptr_inc[2]), .D(n620), .E(
        n619), .F(temp[2]), .Y(n1644) );
  AO222X1 U1886 ( .A(dpl_current[0]), .B(n621), .C(dptr_inc[0]), .D(n620), .E(
        n619), .F(temp[0]), .Y(n1642) );
  MUX4X1 U1887 ( .D0(rn_reg[92]), .D1(rn_reg[84]), .D2(rn_reg[76]), .D3(
        rn_reg[68]), .S0(n372), .S1(n379), .Y(n331) );
  MUX4X1 U1888 ( .D0(rn_reg[220]), .D1(rn_reg[212]), .D2(rn_reg[204]), .D3(
        rn_reg[196]), .S0(n372), .S1(n379), .Y(n336) );
  MUX4X1 U1889 ( .D0(rn_reg[91]), .D1(rn_reg[83]), .D2(rn_reg[75]), .D3(
        rn_reg[67]), .S0(n371), .S1(n378), .Y(n321) );
  MUX4X1 U1890 ( .D0(rn_reg[219]), .D1(rn_reg[211]), .D2(rn_reg[203]), .D3(
        rn_reg[195]), .S0(n371), .S1(n378), .Y(n326) );
  MUX4X1 U1891 ( .D0(rn_reg[60]), .D1(rn_reg[52]), .D2(rn_reg[44]), .D3(
        rn_reg[36]), .S0(n371), .S1(n378), .Y(n330) );
  MUX4X1 U1892 ( .D0(rn_reg[188]), .D1(rn_reg[180]), .D2(rn_reg[172]), .D3(
        rn_reg[164]), .S0(n372), .S1(n379), .Y(n335) );
  MUX4X1 U1893 ( .D0(rn_reg[59]), .D1(rn_reg[51]), .D2(rn_reg[43]), .D3(
        rn_reg[35]), .S0(n371), .S1(n378), .Y(n320) );
  MUX4X1 U1894 ( .D0(rn_reg[187]), .D1(rn_reg[179]), .D2(rn_reg[171]), .D3(
        rn_reg[163]), .S0(n371), .S1(n378), .Y(n325) );
  MUX4X1 U1895 ( .D0(rn_reg[124]), .D1(rn_reg[116]), .D2(rn_reg[108]), .D3(
        rn_reg[100]), .S0(n372), .S1(n379), .Y(n332) );
  MUX4X1 U1896 ( .D0(rn_reg[252]), .D1(rn_reg[244]), .D2(rn_reg[236]), .D3(
        rn_reg[228]), .S0(n372), .S1(n379), .Y(n337) );
  MUX4X1 U1897 ( .D0(rn_reg[123]), .D1(rn_reg[115]), .D2(rn_reg[107]), .D3(
        rn_reg[99]), .S0(n371), .S1(n378), .Y(n322) );
  MUX4X1 U1898 ( .D0(rn_reg[251]), .D1(rn_reg[243]), .D2(rn_reg[235]), .D3(
        rn_reg[227]), .S0(n371), .S1(n378), .Y(n327) );
  MUX4X1 U1899 ( .D0(rn_reg[28]), .D1(rn_reg[20]), .D2(rn_reg[12]), .D3(
        rn_reg[4]), .S0(n371), .S1(n378), .Y(n329) );
  MUX4X1 U1900 ( .D0(rn_reg[156]), .D1(rn_reg[148]), .D2(rn_reg[140]), .D3(
        rn_reg[132]), .S0(n372), .S1(n379), .Y(n334) );
  MUX4X1 U1901 ( .D0(rn_reg[27]), .D1(rn_reg[19]), .D2(rn_reg[11]), .D3(
        rn_reg[3]), .S0(n371), .S1(n378), .Y(n319) );
  MUX4X1 U1902 ( .D0(rn_reg[155]), .D1(rn_reg[147]), .D2(rn_reg[139]), .D3(
        rn_reg[131]), .S0(n371), .S1(n378), .Y(n324) );
  MUX2X1 U1903 ( .D0(n820), .D1(n819), .S(codefetch_s), .Y(n840) );
  NAND21X1 U1904 ( .B(n880), .A(mempsrd), .Y(n820) );
  NAND21X1 U1905 ( .B(stop_r), .A(n725), .Y(n819) );
  AOI211X1 U1906 ( .C(n432), .D(n749), .A(n882), .B(n883), .Y(n880) );
  MUX2X1 U1907 ( .D0(memaddr[0]), .D1(n1642), .S(n622), .Y(N12841) );
  AO21X1 U1908 ( .B(n946), .C(n121), .A(n1034), .Y(n1763) );
  OAI31XL U1909 ( .A(n2017), .B(n1035), .C(n1036), .D(n2166), .Y(n1034) );
  INVX1 U1910 ( .A(israccess), .Y(n2166) );
  NAND21X1 U1911 ( .B(n1037), .A(n1989), .Y(n1036) );
  INVX1 U1912 ( .A(n2189), .Y(n1955) );
  AND2X1 U1913 ( .A(n1747), .B(n2194), .Y(N353) );
  INVX1 U1914 ( .A(ramdatao[3]), .Y(n2128) );
  ENOX1 U1915 ( .A(n2120), .B(n91), .C(N11840), .D(n1275), .Y(dpl_current[2])
         );
  MUX2X1 U1916 ( .D0(n274), .D1(n273), .S(n119), .Y(N11840) );
  MUX4X1 U1917 ( .D0(dpl_reg[2]), .D1(dpl_reg[10]), .D2(dpl_reg[18]), .D3(
        dpl_reg[26]), .S0(n285), .S1(n287), .Y(n274) );
  MUX4X1 U1918 ( .D0(dpl_reg[34]), .D1(dpl_reg[42]), .D2(dpl_reg[50]), .D3(
        dpl_reg[58]), .S0(n285), .S1(n287), .Y(n273) );
  INVX1 U1919 ( .A(temp2_comb[2]), .Y(n2162) );
  INVX1 U1920 ( .A(ramsfraddr[5]), .Y(n1963) );
  INVX1 U1921 ( .A(temp2_comb[1]), .Y(n2126) );
  INVX1 U1922 ( .A(ramsfraddr[6]), .Y(n1962) );
  NOR2X1 U1923 ( .A(n2193), .B(n1683), .Y(n1736) );
  NAND2X1 U1924 ( .A(dps[3]), .B(n1340), .Y(n1336) );
  INVX1 U1925 ( .A(n1396), .Y(n673) );
  NAND41X1 U1926 ( .D(n1390), .A(n1389), .B(n1518), .C(n1388), .Y(n1396) );
  AOI222XL U1927 ( .A(N1763), .B(n1423), .C(temp2_comb[2]), .D(n1909), .E(
        pc_i[10]), .F(n1905), .Y(n1518) );
  AO21X1 U1928 ( .B(n1334), .C(n1572), .A(n1330), .Y(n1389) );
  NAND21X1 U1929 ( .B(n2188), .A(n1955), .Y(n2089) );
  AO222X1 U1930 ( .A(n619), .B(temp[6]), .C(dptr_inc[6]), .D(n620), .E(n621), 
        .F(dpl_current[6]), .Y(n1656) );
  AO222X1 U1931 ( .A(dpl_current[5]), .B(n621), .C(dptr_inc[5]), .D(n620), .E(
        n619), .F(temp[5]), .Y(n1655) );
  AND4X1 U1932 ( .A(n930), .B(n1727), .C(n658), .D(n1499), .Y(n1703) );
  AOI21X1 U1933 ( .B(phase[0]), .C(n1728), .A(n1729), .Y(n1727) );
  NAND2X1 U1934 ( .A(n1726), .B(n2043), .Y(n1728) );
  MUX4X1 U1935 ( .D0(rn_reg[89]), .D1(rn_reg[81]), .D2(rn_reg[73]), .D3(
        rn_reg[65]), .S0(N352), .S1(n376), .Y(n301) );
  MUX4X1 U1936 ( .D0(rn_reg[217]), .D1(rn_reg[209]), .D2(rn_reg[201]), .D3(
        rn_reg[193]), .S0(instr[0]), .S1(n377), .Y(n306) );
  MUX4X1 U1937 ( .D0(rn_reg[93]), .D1(rn_reg[85]), .D2(rn_reg[77]), .D3(
        rn_reg[69]), .S0(n372), .S1(n379), .Y(n341) );
  MUX4X1 U1938 ( .D0(rn_reg[221]), .D1(rn_reg[213]), .D2(rn_reg[205]), .D3(
        rn_reg[197]), .S0(n373), .S1(n380), .Y(n346) );
  MUX4X1 U1939 ( .D0(rn_reg[94]), .D1(rn_reg[86]), .D2(rn_reg[78]), .D3(
        rn_reg[70]), .S0(n373), .S1(n380), .Y(n351) );
  MUX4X1 U1940 ( .D0(rn_reg[222]), .D1(rn_reg[214]), .D2(rn_reg[206]), .D3(
        rn_reg[198]), .S0(n374), .S1(n381), .Y(n356) );
  MUX4X1 U1941 ( .D0(rn_reg[216]), .D1(rn_reg[208]), .D2(rn_reg[200]), .D3(
        rn_reg[192]), .S0(N352), .S1(n376), .Y(n296) );
  MUX4X1 U1942 ( .D0(rn_reg[88]), .D1(rn_reg[80]), .D2(rn_reg[72]), .D3(
        rn_reg[64]), .S0(n370), .S1(N353), .Y(n291) );
  MUX4X1 U1943 ( .D0(rn_reg[57]), .D1(rn_reg[49]), .D2(rn_reg[41]), .D3(
        rn_reg[33]), .S0(n444), .S1(n376), .Y(n300) );
  MUX4X1 U1944 ( .D0(rn_reg[185]), .D1(rn_reg[177]), .D2(rn_reg[169]), .D3(
        rn_reg[161]), .S0(n444), .S1(n376), .Y(n305) );
  MUX4X1 U1945 ( .D0(rn_reg[61]), .D1(rn_reg[53]), .D2(rn_reg[45]), .D3(
        rn_reg[37]), .S0(n372), .S1(n379), .Y(n340) );
  MUX4X1 U1946 ( .D0(rn_reg[189]), .D1(rn_reg[181]), .D2(rn_reg[173]), .D3(
        rn_reg[165]), .S0(n373), .S1(n380), .Y(n345) );
  MUX4X1 U1947 ( .D0(rn_reg[62]), .D1(rn_reg[54]), .D2(rn_reg[46]), .D3(
        rn_reg[38]), .S0(n373), .S1(n380), .Y(n350) );
  MUX4X1 U1948 ( .D0(rn_reg[190]), .D1(rn_reg[182]), .D2(rn_reg[174]), .D3(
        rn_reg[166]), .S0(n373), .S1(n380), .Y(n355) );
  MUX4X1 U1949 ( .D0(rn_reg[184]), .D1(rn_reg[176]), .D2(rn_reg[168]), .D3(
        rn_reg[160]), .S0(N352), .S1(n376), .Y(n295) );
  MUX4X1 U1950 ( .D0(rn_reg[56]), .D1(rn_reg[48]), .D2(rn_reg[40]), .D3(
        rn_reg[32]), .S0(n370), .S1(N353), .Y(n290) );
  MUX4X1 U1951 ( .D0(rn_reg[121]), .D1(rn_reg[113]), .D2(rn_reg[105]), .D3(
        rn_reg[97]), .S0(n444), .S1(n376), .Y(n302) );
  MUX4X1 U1952 ( .D0(rn_reg[249]), .D1(rn_reg[241]), .D2(rn_reg[233]), .D3(
        rn_reg[225]), .S0(n370), .S1(n377), .Y(n307) );
  MUX4X1 U1953 ( .D0(rn_reg[125]), .D1(rn_reg[117]), .D2(rn_reg[109]), .D3(
        rn_reg[101]), .S0(n372), .S1(n379), .Y(n342) );
  MUX4X1 U1954 ( .D0(rn_reg[253]), .D1(rn_reg[245]), .D2(rn_reg[237]), .D3(
        rn_reg[229]), .S0(n373), .S1(n380), .Y(n347) );
  MUX4X1 U1955 ( .D0(rn_reg[126]), .D1(rn_reg[118]), .D2(rn_reg[110]), .D3(
        rn_reg[102]), .S0(n373), .S1(n380), .Y(n352) );
  MUX4X1 U1956 ( .D0(rn_reg[254]), .D1(rn_reg[246]), .D2(rn_reg[238]), .D3(
        rn_reg[230]), .S0(n374), .S1(n381), .Y(n357) );
  MUX4X1 U1957 ( .D0(rn_reg[248]), .D1(rn_reg[240]), .D2(rn_reg[232]), .D3(
        rn_reg[224]), .S0(N352), .S1(n376), .Y(n297) );
  MUX4X1 U1958 ( .D0(rn_reg[120]), .D1(rn_reg[112]), .D2(rn_reg[104]), .D3(
        rn_reg[96]), .S0(n370), .S1(N353), .Y(n292) );
  MUX4X1 U1959 ( .D0(dpl_reg[35]), .D1(dpl_reg[43]), .D2(dpl_reg[51]), .D3(
        dpl_reg[59]), .S0(n286), .S1(n288), .Y(n275) );
  MUX4X1 U1960 ( .D0(dpl_reg[36]), .D1(dpl_reg[44]), .D2(dpl_reg[52]), .D3(
        dpl_reg[60]), .S0(n286), .S1(n288), .Y(n277) );
  MUX4X1 U1961 ( .D0(rn_reg[25]), .D1(rn_reg[17]), .D2(rn_reg[9]), .D3(
        rn_reg[1]), .S0(N352), .S1(n376), .Y(n299) );
  MUX4X1 U1962 ( .D0(rn_reg[153]), .D1(rn_reg[145]), .D2(rn_reg[137]), .D3(
        rn_reg[129]), .S0(N352), .S1(n376), .Y(n304) );
  MUX4X1 U1963 ( .D0(rn_reg[29]), .D1(rn_reg[21]), .D2(rn_reg[13]), .D3(
        rn_reg[5]), .S0(n372), .S1(n379), .Y(n339) );
  MUX4X1 U1964 ( .D0(rn_reg[157]), .D1(rn_reg[149]), .D2(rn_reg[141]), .D3(
        rn_reg[133]), .S0(n373), .S1(n380), .Y(n344) );
  MUX4X1 U1965 ( .D0(rn_reg[30]), .D1(rn_reg[22]), .D2(rn_reg[14]), .D3(
        rn_reg[6]), .S0(n373), .S1(n380), .Y(n349) );
  MUX4X1 U1966 ( .D0(rn_reg[158]), .D1(rn_reg[150]), .D2(rn_reg[142]), .D3(
        rn_reg[134]), .S0(n373), .S1(n380), .Y(n354) );
  MUX4X1 U1967 ( .D0(rn_reg[152]), .D1(rn_reg[144]), .D2(rn_reg[136]), .D3(
        rn_reg[128]), .S0(N352), .S1(n376), .Y(n294) );
  MUX4X1 U1968 ( .D0(rn_reg[24]), .D1(rn_reg[16]), .D2(rn_reg[8]), .D3(
        rn_reg[0]), .S0(n370), .S1(N353), .Y(n289) );
  NAND21X1 U1969 ( .B(n1157), .A(phase[0]), .Y(n739) );
  NAND32X1 U1970 ( .B(n589), .C(n588), .A(n587), .Y(n968) );
  OA22X1 U1971 ( .A(n92), .B(n2141), .C(n2154), .D(n1183), .Y(n587) );
  AO21X1 U1972 ( .B(n1926), .C(acc[7]), .A(n1462), .Y(n589) );
  AO2222XL U1973 ( .A(n2159), .B(n1917), .C(adder_out[5]), .D(n607), .E(acc[4]), .F(n590), .G(n1919), .H(acc[1]), .Y(n588) );
  NAND42X1 U1974 ( .C(n1423), .D(n1611), .A(n1456), .B(n1732), .Y(n1729) );
  AOI21X1 U1975 ( .B(n1733), .C(phase[1]), .A(n1602), .Y(n1732) );
  INVX1 U1976 ( .A(n2034), .Y(n1733) );
  INVX1 U1977 ( .A(n2194), .Y(n1958) );
  NOR2X1 U1978 ( .A(n2105), .B(instr[6]), .Y(n1682) );
  NOR21XL U1979 ( .B(n457), .A(n996), .Y(N515) );
  NOR21XL U1980 ( .B(n757), .A(n995), .Y(n996) );
  OAI21X1 U1981 ( .B(stop), .C(stop_r), .A(n1841), .Y(n757) );
  INVX1 U1982 ( .A(n2188), .Y(n2105) );
  AND2X1 U1983 ( .A(n1670), .B(phase[0]), .Y(n1602) );
  NAND32X1 U1984 ( .B(n586), .C(n585), .A(n584), .Y(n967) );
  OA22X1 U1985 ( .A(n2134), .B(n92), .C(n1967), .D(n1183), .Y(n584) );
  AO21X1 U1986 ( .B(acc[6]), .C(n1926), .A(n1486), .Y(n586) );
  AO2222XL U1987 ( .A(n2140), .B(n1917), .C(adder_out[4]), .D(n607), .E(n590), 
        .F(acc[3]), .G(n1919), .H(acc[0]), .Y(n585) );
  NOR2X1 U1988 ( .A(n442), .B(n2194), .Y(n1117) );
  XNOR2XL U1989 ( .A(acc[4]), .B(n1370), .Y(N11545) );
  INVX1 U1990 ( .A(ramdatao[0]), .Y(n2053) );
  ENOX1 U1991 ( .A(n1709), .B(n2053), .C(sp[0]), .D(n1709), .Y(N12769) );
  INVX1 U1992 ( .A(n600), .Y(dpl_current[3]) );
  MUX2BXL U1993 ( .D0(n2128), .D1(N11839), .S(n1275), .Y(n600) );
  MUX2X1 U1994 ( .D0(n276), .D1(n275), .S(n118), .Y(N11839) );
  MUX4X1 U1995 ( .D0(dpl_reg[3]), .D1(dpl_reg[11]), .D2(dpl_reg[19]), .D3(
        dpl_reg[27]), .S0(n286), .S1(n288), .Y(n276) );
  NOR2X1 U1996 ( .A(n1958), .B(n104), .Y(n903) );
  INVX1 U1997 ( .A(acc[7]), .Y(n1966) );
  ENOX1 U1998 ( .A(n1709), .B(n2064), .C(sp[1]), .D(n1709), .Y(N12770) );
  AO22X1 U1999 ( .A(n394), .B(n1505), .C(pc_ini[14]), .D(n460), .Y(N494) );
  AO22X1 U2000 ( .A(n393), .B(n1504), .C(pc_ini[13]), .D(n460), .Y(N493) );
  AO22X1 U2001 ( .A(n393), .B(n1503), .C(pc_ini[12]), .D(n460), .Y(N492) );
  AO22X1 U2002 ( .A(n393), .B(n1502), .C(pc_ini[11]), .D(n460), .Y(N491) );
  AO22X1 U2003 ( .A(n393), .B(n1506), .C(pc_ini[15]), .D(n460), .Y(N495) );
  NAND3X1 U2004 ( .A(n1731), .B(interrupt), .C(n933), .Y(n930) );
  NOR2X1 U2005 ( .A(n2123), .B(waitcnt[2]), .Y(n1812) );
  NOR2X1 U2006 ( .A(n2138), .B(waitcnt[2]), .Y(n1809) );
  NOR3XL U2007 ( .A(n2042), .B(n2193), .C(n2087), .Y(n932) );
  INVX1 U2008 ( .A(temp2_comb[3]), .Y(n2153) );
  INVX1 U2009 ( .A(n599), .Y(dpl_current[4]) );
  MUX2BXL U2010 ( .D0(n2134), .D1(N11838), .S(n91), .Y(n599) );
  MUX2X1 U2011 ( .D0(n278), .D1(n277), .S(n119), .Y(N11838) );
  MUX4X1 U2012 ( .D0(dpl_reg[4]), .D1(dpl_reg[12]), .D2(dpl_reg[20]), .D3(
        dpl_reg[28]), .S0(n286), .S1(n288), .Y(n278) );
  INVX1 U2013 ( .A(n714), .Y(n1035) );
  AO2222XL U2014 ( .A(temp[7]), .B(n713), .C(n166), .D(n712), .E(n2010), .F(
        n711), .G(ramsfraddr[7]), .H(n710), .Y(n714) );
  INVX1 U2015 ( .A(n1702), .Y(n711) );
  INVX1 U2016 ( .A(n1703), .Y(n712) );
  AOI21BBXL U2017 ( .B(n1374), .C(n1375), .A(n2110), .Y(n1373) );
  AOI211X1 U2018 ( .C(acc[7]), .D(n1376), .A(c), .B(n1377), .Y(n1374) );
  NAND2X1 U2019 ( .A(n1556), .B(n2159), .Y(n1376) );
  NOR43XL U2020 ( .B(n1378), .C(acc[4]), .D(acc[7]), .A(n2154), .Y(n1377) );
  INVX1 U2021 ( .A(n2190), .Y(n448) );
  INVX1 U2022 ( .A(n2190), .Y(n449) );
  INVX1 U2023 ( .A(dps[0]), .Y(n438) );
  INVX1 U2024 ( .A(N352), .Y(n445) );
  NAND3X1 U2025 ( .A(n121), .B(n1957), .C(n932), .Y(n1157) );
  INVX1 U2026 ( .A(N350), .Y(n440) );
  INVX1 U2027 ( .A(ckcon[6]), .Y(n2138) );
  INVX1 U2028 ( .A(n464), .Y(n1690) );
  OAI211X1 U2029 ( .C(n1813), .D(n1812), .A(n1814), .B(n468), .Y(n464) );
  OAI22X1 U2030 ( .A(waitcnt[0]), .B(n2125), .C(waitcnt[1]), .D(n2124), .Y(
        n1813) );
  AOI32X1 U2031 ( .A(n2122), .B(n2124), .C(waitcnt[1]), .D(waitcnt[2]), .E(
        n2123), .Y(n1814) );
  OAI22X1 U2032 ( .A(waitcnt[0]), .B(n2135), .C(waitcnt[1]), .D(n2142), .Y(
        n1810) );
  AOI32X1 U2033 ( .A(n2137), .B(n2142), .C(waitcnt[1]), .D(waitcnt[2]), .E(
        n2138), .Y(n1811) );
  MUX2X1 U2034 ( .D0(n1917), .D1(n546), .S(acc[0]), .Y(n547) );
  AO21X1 U2035 ( .B(n1921), .C(n1225), .A(n2045), .Y(n546) );
  AOI32X1 U2036 ( .A(n2074), .B(n2075), .C(ramdatao[2]), .D(n1338), .E(rs[1]), 
        .Y(n1341) );
  AO222X1 U2037 ( .A(dpl_current[7]), .B(n621), .C(dptr_inc[7]), .D(n620), .E(
        n619), .F(temp[7]), .Y(n1659) );
  MUX4X1 U2038 ( .D0(n367), .D1(n365), .D2(n366), .D3(n364), .S0(n2065), .S1(
        n100), .Y(n368) );
  MUX4X1 U2039 ( .D0(rn_reg[223]), .D1(rn_reg[215]), .D2(rn_reg[207]), .D3(
        rn_reg[199]), .S0(n374), .S1(n381), .Y(n366) );
  MUX4X1 U2040 ( .D0(rn_reg[159]), .D1(rn_reg[151]), .D2(rn_reg[143]), .D3(
        rn_reg[135]), .S0(n374), .S1(n381), .Y(n364) );
  MUX4X1 U2041 ( .D0(rn_reg[255]), .D1(rn_reg[247]), .D2(rn_reg[239]), .D3(
        rn_reg[231]), .S0(n374), .S1(n381), .Y(n367) );
  MUX4X1 U2042 ( .D0(dph_reg[7]), .D1(dph_reg[15]), .D2(dph_reg[23]), .D3(
        dph_reg[31]), .S0(n250), .S1(n246), .Y(n217) );
  MUX4X1 U2043 ( .D0(dpl_reg[7]), .D1(dpl_reg[15]), .D2(dpl_reg[23]), .D3(
        dpl_reg[31]), .S0(n249), .S1(dps[1]), .Y(n201) );
  MUX4X1 U2044 ( .D0(rn_reg[90]), .D1(rn_reg[82]), .D2(rn_reg[74]), .D3(
        rn_reg[66]), .S0(instr[0]), .S1(n377), .Y(n311) );
  MUX4X1 U2045 ( .D0(rn_reg[218]), .D1(rn_reg[210]), .D2(rn_reg[202]), .D3(
        rn_reg[194]), .S0(N352), .S1(n377), .Y(n316) );
  MUX4X1 U2046 ( .D0(rn_reg[95]), .D1(rn_reg[87]), .D2(rn_reg[79]), .D3(
        rn_reg[71]), .S0(n374), .S1(n381), .Y(n361) );
  MUX4X1 U2047 ( .D0(rn_reg[58]), .D1(rn_reg[50]), .D2(rn_reg[42]), .D3(
        rn_reg[34]), .S0(instr[0]), .S1(n377), .Y(n310) );
  MUX4X1 U2048 ( .D0(rn_reg[186]), .D1(rn_reg[178]), .D2(rn_reg[170]), .D3(
        rn_reg[162]), .S0(instr[0]), .S1(n377), .Y(n315) );
  MUX4X1 U2049 ( .D0(rn_reg[191]), .D1(rn_reg[183]), .D2(rn_reg[175]), .D3(
        rn_reg[167]), .S0(n374), .S1(n381), .Y(n365) );
  MUX4X1 U2050 ( .D0(rn_reg[63]), .D1(rn_reg[55]), .D2(rn_reg[47]), .D3(
        rn_reg[39]), .S0(n374), .S1(n381), .Y(n360) );
  MUX4X1 U2051 ( .D0(rn_reg[122]), .D1(rn_reg[114]), .D2(rn_reg[106]), .D3(
        rn_reg[98]), .S0(instr[0]), .S1(n377), .Y(n312) );
  MUX4X1 U2052 ( .D0(rn_reg[250]), .D1(rn_reg[242]), .D2(rn_reg[234]), .D3(
        rn_reg[226]), .S0(instr[0]), .S1(n377), .Y(n317) );
  MUX4X1 U2053 ( .D0(rn_reg[127]), .D1(rn_reg[119]), .D2(rn_reg[111]), .D3(
        rn_reg[103]), .S0(n374), .S1(n381), .Y(n362) );
  MUX4X1 U2054 ( .D0(dpl_reg[38]), .D1(dpl_reg[46]), .D2(dpl_reg[54]), .D3(
        dpl_reg[62]), .S0(n286), .S1(n288), .Y(n281) );
  MUX2X1 U2055 ( .D0(n237), .D1(n236), .S(n245), .Y(dpc[3]) );
  MUX4X1 U2056 ( .D0(dpc_tab[3]), .D1(dpc_tab[9]), .D2(dpc_tab[15]), .D3(
        dpc_tab[21]), .S0(n252), .S1(n248), .Y(n237) );
  MUX4X1 U2057 ( .D0(dpc_tab[27]), .D1(dpc_tab[33]), .D2(dpc_tab[39]), .D3(
        dpc_tab[45]), .S0(n252), .S1(n248), .Y(n236) );
  MUX2X1 U2058 ( .D0(n241), .D1(n240), .S(n245), .Y(dpc[1]) );
  MUX4X1 U2059 ( .D0(dpc_tab[1]), .D1(dpc_tab[7]), .D2(dpc_tab[13]), .D3(
        dpc_tab[19]), .S0(n252), .S1(n248), .Y(n241) );
  MUX4X1 U2060 ( .D0(dpc_tab[25]), .D1(dpc_tab[31]), .D2(dpc_tab[37]), .D3(
        dpc_tab[43]), .S0(n252), .S1(n248), .Y(n240) );
  MUX4X1 U2061 ( .D0(dph_reg[39]), .D1(dph_reg[47]), .D2(dph_reg[55]), .D3(
        dph_reg[63]), .S0(n250), .S1(n246), .Y(n216) );
  MUX4X1 U2062 ( .D0(dpl_reg[38]), .D1(dpl_reg[46]), .D2(dpl_reg[54]), .D3(
        dpl_reg[62]), .S0(n249), .S1(dps[1]), .Y(n202) );
  MUX4X1 U2063 ( .D0(dpl_reg[39]), .D1(dpl_reg[47]), .D2(dpl_reg[55]), .D3(
        dpl_reg[63]), .S0(n249), .S1(dps[1]), .Y(n200) );
  MUX4X1 U2064 ( .D0(rn_reg[26]), .D1(rn_reg[18]), .D2(rn_reg[10]), .D3(
        rn_reg[2]), .S0(n444), .S1(n377), .Y(n309) );
  MUX4X1 U2065 ( .D0(rn_reg[154]), .D1(rn_reg[146]), .D2(rn_reg[138]), .D3(
        rn_reg[130]), .S0(N352), .S1(n377), .Y(n314) );
  MUX4X1 U2066 ( .D0(rn_reg[31]), .D1(rn_reg[23]), .D2(rn_reg[15]), .D3(
        rn_reg[7]), .S0(n374), .S1(n381), .Y(n359) );
  MUX2BXL U2067 ( .D0(n190), .D1(ramdatao[7]), .S(n580), .Y(n1566) );
  MUX2IX1 U2068 ( .D0(n368), .D1(n363), .S(n2066), .Y(n190) );
  OR2X1 U2069 ( .A(ramsfraddr[3]), .B(ramsfraddr[4]), .Y(n509) );
  INVX1 U2070 ( .A(n104), .Y(n1957) );
  INVX1 U2071 ( .A(n2191), .Y(n1956) );
  OR2X1 U2072 ( .A(memrd), .B(memwr), .Y(n468) );
  AO222X1 U2073 ( .A(n11), .B(pc_o[5]), .C(n13), .D(n1483), .E(pc_ini[5]), .F(
        n462), .Y(N485) );
  AO222X1 U2074 ( .A(n12), .B(memaddr[6]), .C(n14), .D(n1484), .E(pc_ini[6]), 
        .F(n461), .Y(N486) );
  AO222X1 U2075 ( .A(n11), .B(N1761), .C(n13), .D(n1476), .E(pc_ini[0]), .F(
        n462), .Y(N480) );
  AO222X1 U2076 ( .A(n12), .B(n2185), .C(n14), .D(n1485), .E(pc_ini[7]), .F(
        n459), .Y(N487) );
  AO222X1 U2077 ( .A(n11), .B(pc_o[4]), .C(n13), .D(n1481), .E(pc_ini[4]), .F(
        n460), .Y(N484) );
  AO222X1 U2078 ( .A(n12), .B(memaddr[3]), .C(n14), .D(n1479), .E(pc_ini[3]), 
        .F(n460), .Y(N483) );
  AO222X1 U2079 ( .A(n11), .B(pc_o[2]), .C(n13), .D(n1478), .E(pc_ini[2]), .F(
        n462), .Y(N482) );
  AO222X1 U2080 ( .A(n12), .B(memaddr[10]), .C(n14), .D(n1501), .E(pc_ini[10]), 
        .F(n458), .Y(N490) );
  AO222X1 U2081 ( .A(n11), .B(pc_o[9]), .C(n13), .D(n1500), .E(pc_ini[9]), .F(
        n458), .Y(N489) );
  AO222X1 U2082 ( .A(n12), .B(memaddr[8]), .C(n14), .D(n1491), .E(pc_ini[8]), 
        .F(n458), .Y(N488) );
  AO222X1 U2083 ( .A(n11), .B(memaddr[1]), .C(n13), .D(n1477), .E(pc_ini[1]), 
        .F(n459), .Y(N481) );
  OAI21X1 U2084 ( .B(dec_accop[7]), .C(n1381), .A(n115), .Y(n1658) );
  AOI22X1 U2085 ( .A(n2067), .B(ramdatao[4]), .C(n1168), .D(rs[1]), .Y(n1188)
         );
  OR2X1 U2086 ( .A(mempswr), .B(mempsrd), .Y(n470) );
  INVX1 U2087 ( .A(n535), .Y(n580) );
  NAND41X1 U2088 ( .D(n8), .A(n1743), .B(n1741), .C(n1742), .Y(n535) );
  XNOR2XL U2089 ( .A(n2066), .B(ramsfraddr[4]), .Y(n1741) );
  XNOR2XL U2090 ( .A(n2065), .B(ramsfraddr[3]), .Y(n1742) );
  INVX1 U2091 ( .A(n2193), .Y(n2106) );
  EORX1 U2092 ( .A(phase[1]), .B(n908), .C(n1738), .D(n123), .Y(n1713) );
  OAI31XL U2093 ( .A(n1739), .B(n1952), .C(n2080), .D(n104), .Y(n1738) );
  OAI21X1 U2094 ( .B(n1955), .C(n960), .A(n2087), .Y(n1739) );
  AND2X1 U2095 ( .A(dec_accop[14]), .B(n115), .Y(n1360) );
  MUX2X1 U2096 ( .D0(n604), .D1(n1550), .S(acc[1]), .Y(n526) );
  AOI21X1 U2097 ( .B(n80), .C(n2126), .A(n2045), .Y(n1550) );
  MUX2X1 U2098 ( .D0(n604), .D1(n1532), .S(acc[2]), .Y(n559) );
  AOI21X1 U2099 ( .B(n80), .C(n2162), .A(n2045), .Y(n1532) );
  AO21X1 U2100 ( .B(n2184), .C(n982), .A(n462), .Y(N520) );
  MUX2X1 U2101 ( .D0(p2sel), .D1(n1401), .S(n981), .Y(n982) );
  INVX1 U2102 ( .A(n598), .Y(dpl_current[6]) );
  MUX2BXL U2103 ( .D0(n2136), .D1(N11836), .S(n1275), .Y(n598) );
  MUX2X1 U2104 ( .D0(n282), .D1(n281), .S(n119), .Y(N11836) );
  MUX4X1 U2105 ( .D0(dpl_reg[6]), .D1(dpl_reg[14]), .D2(dpl_reg[22]), .D3(
        dpl_reg[30]), .S0(n286), .S1(n288), .Y(n282) );
  NAND2X1 U2106 ( .A(dec_accop[0]), .B(n116), .Y(n1226) );
  NOR2X1 U2107 ( .A(n2193), .B(n104), .Y(n1124) );
  NAND2X1 U2108 ( .A(n1594), .B(instr[4]), .Y(n1821) );
  MUX2BXL U2109 ( .D0(n2044), .D1(n1366), .S(acc[0]), .Y(n542) );
  ENOX1 U2110 ( .A(n1709), .B(n2120), .C(sp[2]), .D(n1709), .Y(N12771) );
  ENOX1 U2111 ( .A(n1709), .B(n2128), .C(sp[3]), .D(n1709), .Y(N12772) );
  ENOX1 U2112 ( .A(n107), .B(n2134), .C(sp[4]), .D(n1709), .Y(N12773) );
  NOR2X1 U2113 ( .A(n2106), .B(instr[4]), .Y(n901) );
  NOR2X1 U2114 ( .A(n429), .B(n104), .Y(n933) );
  INVX1 U2115 ( .A(acc[3]), .Y(n2154) );
  INVX1 U2116 ( .A(acc[5]), .Y(n2159) );
  ENOX1 U2117 ( .A(n2141), .B(n91), .C(N11837), .D(n1275), .Y(dpl_current[5])
         );
  MUX2X1 U2118 ( .D0(n280), .D1(n279), .S(n118), .Y(N11837) );
  MUX4X1 U2119 ( .D0(dpl_reg[5]), .D1(dpl_reg[13]), .D2(dpl_reg[21]), .D3(
        dpl_reg[29]), .S0(n286), .S1(n288), .Y(n280) );
  MUX4X1 U2120 ( .D0(dpl_reg[37]), .D1(dpl_reg[45]), .D2(dpl_reg[53]), .D3(
        dpl_reg[61]), .S0(n286), .S1(n288), .Y(n279) );
  NAND2X1 U2121 ( .A(dec_accop[1]), .B(n115), .Y(n1224) );
  NAND2X1 U2122 ( .A(dec_accop[3]), .B(n115), .Y(n1660) );
  INVX1 U2123 ( .A(phase[1]), .Y(n2077) );
  NAND2X1 U2124 ( .A(dec_accop[13]), .B(n116), .Y(n1653) );
  OAI222XL U2125 ( .A(n1463), .B(n2158), .C(n1464), .D(n2159), .E(n2048), .F(
        n1556), .Y(n1462) );
  AOI221XL U2126 ( .A(acc[5]), .B(n1366), .C(n1921), .D(n2159), .E(n2047), .Y(
        n1463) );
  AOI21X1 U2127 ( .B(n1921), .C(n2158), .A(n2045), .Y(n1464) );
  OAI222XL U2128 ( .A(n1487), .B(n2156), .C(n1488), .D(n2140), .E(n2048), .F(
        n2159), .Y(n1486) );
  AOI221XL U2129 ( .A(n1366), .B(acc[4]), .C(n1921), .D(n2140), .E(n2047), .Y(
        n1487) );
  AOI21X1 U2130 ( .B(n1921), .C(n2156), .A(n2045), .Y(n1488) );
  OAI222XL U2131 ( .A(n1436), .B(n2139), .C(n1437), .D(n1556), .E(n2048), .F(
        n1966), .Y(n1435) );
  AOI221XL U2132 ( .A(acc[6]), .B(n1366), .C(n1921), .D(n1556), .E(n2047), .Y(
        n1436) );
  AOI21X1 U2133 ( .B(n1921), .C(n2139), .A(n2045), .Y(n1437) );
  INVX1 U2134 ( .A(temp2_comb[4]), .Y(n2156) );
  AOI211X1 U2135 ( .C(n693), .D(n1804), .A(n459), .B(n1274), .Y(n1290) );
  OAI21X1 U2136 ( .B(temp2_comb[7]), .C(n2044), .A(n1409), .Y(n1408) );
  OAI221XL U2137 ( .A(n2076), .B(n1074), .C(n678), .D(n1065), .E(n457), .Y(
        n1878) );
  INVX1 U2138 ( .A(newinstrlock), .Y(n2076) );
  OAI22AX1 U2139 ( .D(stop), .C(n681), .A(n1960), .B(n678), .Y(n1880) );
  OAI22AX1 U2140 ( .D(idle), .C(n681), .A(n678), .B(n1953), .Y(n1879) );
  OAI21X1 U2141 ( .B(n1406), .C(n2160), .A(n1407), .Y(n1400) );
  AOI221XL U2142 ( .A(n1366), .B(acc[7]), .C(n1921), .D(n1966), .E(n2047), .Y(
        n1406) );
  AOI32X1 U2143 ( .A(n529), .B(n1227), .C(acc[0]), .D(acc[7]), .E(n1408), .Y(
        n1407) );
  NAND3X1 U2144 ( .A(n2119), .B(n2121), .C(ramsfraddr[0]), .Y(n1002) );
  NAND2X1 U2145 ( .A(instr[4]), .B(n2106), .Y(n1689) );
  NOR3XL U2146 ( .A(n1744), .B(n1745), .C(n1746), .Y(n1743) );
  XNOR2XL U2147 ( .A(n442), .B(ramsfraddr[0]), .Y(n1745) );
  XNOR2XL U2148 ( .A(n100), .B(n2121), .Y(n1746) );
  XNOR2XL U2149 ( .A(N353), .B(n2119), .Y(n1744) );
  NAND32X1 U2150 ( .B(n563), .C(n562), .A(n561), .Y(n1361) );
  OAI22X1 U2151 ( .A(n1227), .B(n2120), .C(n2127), .D(n1356), .Y(n563) );
  AOI222XL U2152 ( .A(acc[6]), .B(n1919), .C(n608), .D(acc[3]), .E(
        adder_out[2]), .F(n607), .Y(n561) );
  OAI211X1 U2153 ( .C(n1531), .D(n2162), .A(n559), .B(n558), .Y(n562) );
  INVX1 U2154 ( .A(ckcon[2]), .Y(n2123) );
  INVX1 U2155 ( .A(ckcon[1]), .Y(n2124) );
  INVX1 U2156 ( .A(ckcon[5]), .Y(n2142) );
  INVX1 U2157 ( .A(ckcon[4]), .Y(n2135) );
  INVX1 U2158 ( .A(ckcon[0]), .Y(n2125) );
  AND2X1 U2159 ( .A(dec_accop[2]), .B(n116), .Y(n191) );
  NAND43X1 U2160 ( .B(dec_accop[18]), .C(n1735), .D(n1222), .A(n1927), .Y(
        n1183) );
  MUX2BXL U2161 ( .D0(n2134), .D1(pmw), .S(n686), .Y(n1941) );
  AO222X1 U2162 ( .A(dph_current[1]), .B(n616), .C(dptr_inc[9]), .D(n99), .E(
        n1307), .F(temp[1]), .Y(n1613) );
  AO222X1 U2163 ( .A(dph_current[2]), .B(n616), .C(dptr_inc[10]), .D(n99), .E(
        n1307), .F(temp[2]), .Y(n1615) );
  AO222X1 U2164 ( .A(dph_current[0]), .B(n616), .C(dptr_inc[8]), .D(n620), .E(
        n1307), .F(temp[0]), .Y(n1612) );
  NAND21X1 U2165 ( .B(n1821), .A(n104), .Y(n2081) );
  MUX2X1 U2166 ( .D0(n239), .D1(n238), .S(n245), .Y(dpc[2]) );
  MUX4X1 U2167 ( .D0(dpc_tab[2]), .D1(dpc_tab[8]), .D2(dpc_tab[14]), .D3(
        dpc_tab[20]), .S0(n252), .S1(n248), .Y(n239) );
  MUX4X1 U2168 ( .D0(dpc_tab[26]), .D1(dpc_tab[32]), .D2(dpc_tab[38]), .D3(
        dpc_tab[44]), .S0(n252), .S1(n248), .Y(n238) );
  NAND21X1 U2169 ( .B(n383), .A(dec_accop[15]), .Y(n1657) );
  NOR42XL U2170 ( .C(n1954), .D(n767), .A(phase[5]), .B(n940), .Y(n768) );
  NAND3X1 U2171 ( .A(n429), .B(n2078), .C(n124), .Y(n940) );
  NAND21X1 U2172 ( .B(n383), .A(dec_accop[17]), .Y(n1222) );
  AO21X1 U2173 ( .B(n1573), .C(phase[1]), .A(n651), .Y(n647) );
  NAND21X1 U2174 ( .B(instr[4]), .A(n2194), .Y(n2098) );
  NAND21X1 U2175 ( .B(n383), .A(dec_accop[16]), .Y(n487) );
  NAND32X1 U2176 ( .B(n611), .C(n610), .A(n609), .Y(n868) );
  OAI22X1 U2177 ( .A(n2128), .B(n1227), .C(n1967), .D(n1356), .Y(n611) );
  OAI211X1 U2178 ( .C(n1513), .D(n2153), .A(n606), .B(n605), .Y(n610) );
  AOI222XL U2179 ( .A(n1919), .B(acc[7]), .C(n608), .D(acc[4]), .E(
        adder_out[3]), .F(n607), .Y(n609) );
  OAI211X1 U2180 ( .C(n1384), .D(n2169), .A(n1445), .B(n1446), .Y(n1055) );
  AOI222XL U2181 ( .A(memdatai[5]), .B(n1387), .C(temp2_comb[5]), .D(n1914), 
        .E(n1924), .F(n2012), .Y(n1446) );
  AOI22XL U2182 ( .A(sfrdatai[5]), .B(n1915), .C(n968), .D(n1391), .Y(n1445)
         );
  OAI211X1 U2183 ( .C(n1384), .D(n2168), .A(n1425), .B(n1426), .Y(n1057) );
  AOI222XL U2184 ( .A(memdatai[6]), .B(n1387), .C(temp2_comb[6]), .D(n1914), 
        .E(n1924), .F(n2011), .Y(n1426) );
  AOI22XL U2185 ( .A(sfrdatai[6]), .B(n1915), .C(n969), .D(n1391), .Y(n1425)
         );
  OAI211X1 U2186 ( .C(n1384), .D(n2170), .A(n1465), .B(n1466), .Y(n1056) );
  AOI222XL U2187 ( .A(memdatai[4]), .B(n1387), .C(temp2_comb[4]), .D(n1914), 
        .E(n1924), .F(n2013), .Y(n1466) );
  OAI31XL U2188 ( .A(n1032), .B(n2130), .C(n1941), .D(n1877), .Y(n736) );
  AOI32X1 U2189 ( .A(n2072), .B(n1032), .C(ckcon[7]), .D(n1941), .E(n2069), 
        .Y(n1877) );
  INVX1 U2190 ( .A(n1031), .Y(n2069) );
  NAND21X1 U2191 ( .B(instr[6]), .A(n1331), .Y(n2093) );
  OAI221X1 U2192 ( .A(n1954), .B(n481), .C(n480), .D(n767), .E(n479), .Y(n2019) );
  AND3X1 U2193 ( .A(n1874), .B(n897), .C(n2035), .Y(n481) );
  INVX1 U2194 ( .A(n751), .Y(n480) );
  AOI222XL U2195 ( .A(n1844), .B(phase[1]), .C(n1843), .D(phase[0]), .E(n1842), 
        .F(phase[2]), .Y(n479) );
  NAND21X1 U2196 ( .B(n383), .A(dec_accop[18]), .Y(n1654) );
  MUX2X1 U2197 ( .D0(n243), .D1(n242), .S(n245), .Y(dpc[0]) );
  MUX4X1 U2198 ( .D0(dpc_tab[0]), .D1(dpc_tab[6]), .D2(dpc_tab[12]), .D3(
        dpc_tab[18]), .S0(n252), .S1(n248), .Y(n243) );
  MUX4X1 U2199 ( .D0(dpc_tab[24]), .D1(dpc_tab[30]), .D2(dpc_tab[36]), .D3(
        dpc_tab[42]), .S0(n252), .S1(n248), .Y(n242) );
  OAI211X1 U2200 ( .C(n1467), .D(n1903), .A(n1492), .B(n1493), .Y(n1684) );
  AOI222XL U2201 ( .A(memdatai[3]), .B(n1387), .C(temp2_comb[3]), .D(n1914), 
        .E(n1924), .F(n2014), .Y(n1493) );
  AOI22XL U2202 ( .A(sfrdatai[3]), .B(n1915), .C(ramdatai[3]), .D(n1494), .Y(
        n1492) );
  MUX2X1 U2203 ( .D0(n211), .D1(n210), .S(n244), .Y(dpl[2]) );
  MUX4X1 U2204 ( .D0(dpl_reg[2]), .D1(dpl_reg[10]), .D2(dpl_reg[18]), .D3(
        dpl_reg[26]), .S0(dps[0]), .S1(N350), .Y(n211) );
  MUX4X1 U2205 ( .D0(dpl_reg[34]), .D1(dpl_reg[42]), .D2(dpl_reg[50]), .D3(
        dpl_reg[58]), .S0(dps[0]), .S1(N350), .Y(n210) );
  MUX2X1 U2206 ( .D0(n227), .D1(n226), .S(n245), .Y(dph[2]) );
  MUX4X1 U2207 ( .D0(dph_reg[2]), .D1(dph_reg[10]), .D2(dph_reg[18]), .D3(
        dph_reg[26]), .S0(n251), .S1(n247), .Y(n227) );
  MUX4X1 U2208 ( .D0(dph_reg[34]), .D1(dph_reg[42]), .D2(dph_reg[50]), .D3(
        dph_reg[58]), .S0(n251), .S1(n247), .Y(n226) );
  AOI22X1 U2209 ( .A(ramdatao[3]), .B(n2070), .C(ckcon[3]), .D(n1032), .Y(
        n1031) );
  INVX1 U2210 ( .A(n1383), .Y(n1970) );
  OAI211X1 U2211 ( .C(n1384), .D(n2167), .A(n1385), .B(n1386), .Y(n1383) );
  AOI222XL U2212 ( .A(memdatai[7]), .B(n1387), .C(n1914), .D(temp2_comb[7]), 
        .E(n1924), .F(n2010), .Y(n1386) );
  XNOR2XL U2213 ( .A(acc[6]), .B(n1370), .Y(N11547) );
  XNOR2XL U2214 ( .A(acc[5]), .B(n1370), .Y(N11546) );
  INVX1 U2215 ( .A(ramdatao[1]), .Y(n2064) );
  NOR3XL U2216 ( .A(n2030), .B(n104), .C(n2095), .Y(n1835) );
  MUX2X1 U2217 ( .D0(n604), .D1(n1514), .S(acc[3]), .Y(n606) );
  AOI21X1 U2218 ( .B(n80), .C(n2153), .A(n2045), .Y(n1514) );
  MUX2X1 U2219 ( .D0(n225), .D1(n224), .S(n245), .Y(dph[3]) );
  MUX4X1 U2220 ( .D0(dph_reg[3]), .D1(dph_reg[11]), .D2(dph_reg[19]), .D3(
        dph_reg[27]), .S0(n251), .S1(n247), .Y(n225) );
  MUX4X1 U2221 ( .D0(dph_reg[35]), .D1(dph_reg[43]), .D2(dph_reg[51]), .D3(
        dph_reg[59]), .S0(n251), .S1(n247), .Y(n224) );
  MUX2X1 U2222 ( .D0(n229), .D1(n228), .S(n245), .Y(dph[1]) );
  MUX4X1 U2223 ( .D0(dph_reg[1]), .D1(dph_reg[9]), .D2(dph_reg[17]), .D3(
        dph_reg[25]), .S0(n251), .S1(n247), .Y(n229) );
  MUX4X1 U2224 ( .D0(dph_reg[33]), .D1(dph_reg[41]), .D2(dph_reg[49]), .D3(
        dph_reg[57]), .S0(n251), .S1(n247), .Y(n228) );
  BUFX3 U2225 ( .A(N1761), .Y(pc_o[0]) );
  NOR2X1 U2226 ( .A(n2082), .B(n2188), .Y(n1598) );
  ENOX1 U2227 ( .A(n107), .B(n2141), .C(sp[5]), .D(n107), .Y(N12774) );
  INVX1 U2228 ( .A(ramdatao[2]), .Y(n2120) );
  AND2X1 U2229 ( .A(dec_accop[11]), .B(n116), .Y(n1650) );
  AOI21AX1 U2230 ( .B(n630), .C(n1961), .A(n193), .Y(n192) );
  NAND4X1 U2231 ( .A(n629), .B(phase[1]), .C(n628), .D(n627), .Y(n193) );
  NAND2X1 U2232 ( .A(dec_accop[4]), .B(n116), .Y(n1223) );
  NAND2X1 U2233 ( .A(dec_accop[12]), .B(n116), .Y(n1649) );
  INVX1 U2234 ( .A(ramsfraddr[3]), .Y(n2132) );
  INVX1 U2235 ( .A(interrupt), .Y(n2104) );
  NAND2X1 U2236 ( .A(dec_accop[5]), .B(n115), .Y(n1652) );
  NAND2X1 U2237 ( .A(dec_accop[6]), .B(n115), .Y(n1651) );
  AND2X1 U2238 ( .A(sfroe_r), .B(waitstaten), .Y(sfroe) );
  OAI22X1 U2239 ( .A(n2193), .B(n1866), .C(n2030), .D(n2095), .Y(n895) );
  AOI211X1 U2240 ( .C(n1948), .D(n2105), .A(n1895), .B(n1867), .Y(n1866) );
  AOI21X1 U2241 ( .B(n121), .C(n736), .A(n2105), .Y(n1867) );
  AOI21X1 U2242 ( .B(n627), .C(phase[1]), .A(n623), .Y(n194) );
  NOR2X1 U2243 ( .A(n1957), .B(n121), .Y(n1740) );
  INVX1 U2244 ( .A(temp2_comb[5]), .Y(n2158) );
  NOR2X1 U2245 ( .A(n2132), .B(ramsfraddr[4]), .Y(n1010) );
  OAI22X1 U2246 ( .A(instr[5]), .B(n887), .C(n1862), .D(n1863), .Y(n1842) );
  AOI22X1 U2247 ( .A(n1636), .B(n1117), .C(n890), .D(n891), .Y(n1863) );
  AOI32X1 U2248 ( .A(n901), .B(n63), .C(interrupt), .D(instr[6]), .E(n895), 
        .Y(n1862) );
  AOI221XL U2249 ( .A(acc[3]), .B(n1366), .C(n80), .D(n2154), .E(n2047), .Y(
        n1513) );
  AOI221XL U2250 ( .A(acc[1]), .B(n1366), .C(n1921), .D(n2127), .E(n2047), .Y(
        n1549) );
  AOI221XL U2251 ( .A(acc[2]), .B(n1366), .C(n1921), .D(n1967), .E(n2047), .Y(
        n1531) );
  INVX1 U2252 ( .A(dps[2]), .Y(n441) );
  NAND3X1 U2253 ( .A(ramsfraddr[2]), .B(ramsfraddr[0]), .C(ramsfraddr[1]), .Y(
        n1006) );
  NAND3X1 U2254 ( .A(ramsfraddr[2]), .B(n2071), .C(ramsfraddr[1]), .Y(n1005)
         );
  INVX1 U2255 ( .A(n564), .Y(n1994) );
  OAI211X1 U2256 ( .C(n1467), .D(n1912), .A(n1516), .B(n1517), .Y(n564) );
  AOI222XL U2257 ( .A(memdatai[2]), .B(n1387), .C(temp2_comb[2]), .D(n1914), 
        .E(n1924), .F(n2015), .Y(n1517) );
  AOI22XL U2258 ( .A(sfrdatai[2]), .B(n1915), .C(ramdatai[2]), .D(n1494), .Y(
        n1516) );
  AO222X1 U2259 ( .A(dph_current[3]), .B(n616), .C(dptr_inc[11]), .D(n99), .E(
        n1307), .F(temp[3]), .Y(n1616) );
  AO222X1 U2260 ( .A(dph_current[4]), .B(n616), .C(dptr_inc[12]), .D(n99), .E(
        n1307), .F(temp[4]), .Y(n1617) );
  AO222X1 U2261 ( .A(dph_current[5]), .B(n616), .C(dptr_inc[13]), .D(n99), .E(
        n1307), .F(temp[5]), .Y(n1621) );
  OAI21X1 U2262 ( .B(n431), .C(n507), .A(n1622), .Y(n1387) );
  OAI31XL U2263 ( .A(n1152), .B(n1624), .C(n1625), .D(phase[0]), .Y(n1622) );
  AND3X1 U2264 ( .A(n811), .B(n506), .C(n505), .Y(n507) );
  AND3X1 U2265 ( .A(n1948), .B(n1626), .C(n89), .Y(n1624) );
  MUX2X1 U2266 ( .D0(n1969), .D1(n1968), .S(N345), .Y(N11584) );
  MUX4X1 U2267 ( .D0(temp[0]), .D1(temp[1]), .D2(temp[2]), .D3(temp[3]), .S0(
        N343), .S1(N344), .Y(n1969) );
  MUX4X1 U2268 ( .D0(temp[4]), .D1(temp[5]), .D2(temp[6]), .D3(temp[7]), .S0(
        N343), .S1(N344), .Y(n1968) );
  MUX4X1 U2269 ( .D0(dpl_reg[35]), .D1(dpl_reg[43]), .D2(dpl_reg[51]), .D3(
        dpl_reg[59]), .S0(dps[0]), .S1(N350), .Y(n208) );
  MUX2X1 U2270 ( .D0(n233), .D1(n232), .S(n245), .Y(dpc[5]) );
  MUX4X1 U2271 ( .D0(dpc_tab[5]), .D1(dpc_tab[11]), .D2(dpc_tab[17]), .D3(
        dpc_tab[23]), .S0(n251), .S1(n247), .Y(n233) );
  MUX4X1 U2272 ( .D0(dpc_tab[29]), .D1(dpc_tab[35]), .D2(dpc_tab[41]), .D3(
        dpc_tab[47]), .S0(n251), .S1(n247), .Y(n232) );
  MUX4X1 U2273 ( .D0(dpl_reg[33]), .D1(dpl_reg[41]), .D2(dpl_reg[49]), .D3(
        dpl_reg[57]), .S0(n249), .S1(N350), .Y(n212) );
  MUX2X1 U2274 ( .D0(n235), .D1(n234), .S(n245), .Y(dpc[4]) );
  MUX4X1 U2275 ( .D0(dpc_tab[4]), .D1(dpc_tab[10]), .D2(dpc_tab[16]), .D3(
        dpc_tab[22]), .S0(n252), .S1(n248), .Y(n235) );
  MUX4X1 U2276 ( .D0(dpc_tab[28]), .D1(dpc_tab[34]), .D2(dpc_tab[40]), .D3(
        dpc_tab[46]), .S0(n252), .S1(n248), .Y(n234) );
  AO21X1 U2277 ( .B(N345), .C(n2036), .A(n1480), .Y(n1303) );
  OAI21BBX1 U2278 ( .A(n1344), .B(phase[0]), .C(n195), .Y(n1569) );
  OAI21X1 U2279 ( .B(n978), .C(n977), .A(phase[1]), .Y(n195) );
  AO21X1 U2280 ( .B(n1635), .C(n512), .A(n519), .Y(n537) );
  AOI32X1 U2281 ( .A(n1636), .B(n1116), .C(phase[3]), .D(n432), .E(n1637), .Y(
        n1635) );
  NAND21X1 U2282 ( .B(n511), .A(phase[2]), .Y(n512) );
  NAND21X1 U2283 ( .B(n1625), .A(n1638), .Y(n1637) );
  NAND21X1 U2284 ( .B(n1539), .A(n1589), .Y(n1540) );
  OAI32X1 U2285 ( .A(n430), .B(n1590), .C(n64), .D(n1591), .E(n125), .Y(n1589)
         );
  AOI32X1 U2286 ( .A(n1952), .B(n89), .C(n370), .D(n1594), .E(n903), .Y(n1590)
         );
  AOI22X1 U2287 ( .A(n1892), .B(n1593), .C(n1952), .D(instr[3]), .Y(n1591) );
  AOI22BXL U2288 ( .B(n1601), .A(phase[1]), .D(n1748), .C(phase[0]), .Y(n1716)
         );
  AOI211X1 U2289 ( .C(n1749), .D(n1907), .A(n1750), .B(n1751), .Y(n1748) );
  NOR21XL U2290 ( .B(n960), .A(n1958), .Y(n1749) );
  NAND41X1 U2291 ( .D(n1674), .A(n2034), .B(n1601), .C(n1752), .Y(n1750) );
  NOR2X1 U2292 ( .A(n1955), .B(n2188), .Y(n1839) );
  AO22X1 U2293 ( .A(n750), .B(phase[3]), .C(n748), .D(phase[2]), .Y(n882) );
  ENOX1 U2294 ( .A(n107), .B(n2136), .C(sp[6]), .D(n107), .Y(N12775) );
  AND4X1 U2295 ( .A(n1633), .B(n2081), .C(n2091), .D(n510), .Y(n511) );
  INVX1 U2296 ( .A(n1162), .Y(n510) );
  AOI31X1 U2297 ( .A(n1117), .B(instr[2]), .C(n2080), .D(n909), .Y(n1633) );
  NOR2X1 U2298 ( .A(n2106), .B(n104), .Y(n912) );
  INVX1 U2299 ( .A(phase[2]), .Y(n2078) );
  INVX1 U2300 ( .A(ramdatao[4]), .Y(n2134) );
  ENOX1 U2301 ( .A(n107), .B(n2130), .C(sp[7]), .D(n107), .Y(N12776) );
  ENOX1 U2302 ( .A(n2130), .B(n1275), .C(N11835), .D(n91), .Y(dpl_current[7])
         );
  MUX2X1 U2303 ( .D0(n284), .D1(n283), .S(n118), .Y(N11835) );
  MUX4X1 U2304 ( .D0(dpl_reg[7]), .D1(dpl_reg[15]), .D2(dpl_reg[23]), .D3(
        dpl_reg[31]), .S0(n286), .S1(n288), .Y(n284) );
  MUX4X1 U2305 ( .D0(dpl_reg[39]), .D1(dpl_reg[47]), .D2(dpl_reg[55]), .D3(
        dpl_reg[63]), .S0(n286), .S1(n288), .Y(n283) );
  AOI33X1 U2306 ( .A(n1212), .B(n2133), .C(n1213), .D(c), .E(n2117), .F(n2052), 
        .Y(n1210) );
  INVX1 U2307 ( .A(n1212), .Y(n2052) );
  INVX1 U2308 ( .A(N11584), .Y(n2117) );
  OAI22X1 U2309 ( .A(instr[5]), .B(n887), .C(n888), .D(n889), .Y(n748) );
  AOI21X1 U2310 ( .B(n890), .C(n891), .A(n892), .Y(n889) );
  AOI32X1 U2311 ( .A(n893), .B(n63), .C(n894), .D(instr[6]), .E(n895), .Y(n888) );
  OAI31XL U2312 ( .A(n2104), .B(instr[4]), .C(instr[1]), .D(n896), .Y(n893) );
  NOR3XL U2313 ( .A(n2194), .B(n104), .C(n2097), .Y(n1860) );
  INVX1 U2314 ( .A(temp2_comb[6]), .Y(n2139) );
  NAND2X1 U2315 ( .A(n121), .B(n2194), .Y(n737) );
  AOI22X1 U2316 ( .A(n1205), .B(n1206), .C(dec_cop[0]), .D(n116), .Y(n1204) );
  GEN2XL U2317 ( .D(n2051), .E(c), .C(n1207), .B(N11584), .A(n1208), .Y(n1205)
         );
  INVX1 U2318 ( .A(n1214), .Y(n2051) );
  NOR4XL U2319 ( .A(n1207), .B(n1209), .C(n1210), .D(n1211), .Y(n1208) );
  OAI211X1 U2320 ( .C(instr[5]), .D(n1853), .A(n1854), .B(n1855), .Y(n1843) );
  OAI21BBX1 U2321 ( .A(n16), .B(n1849), .C(instr[3]), .Y(n1854) );
  AOI221XL U2322 ( .A(instr[3]), .B(n57), .C(n1118), .D(n1955), .E(n1861), .Y(
        n1853) );
  AOI22AXL U2323 ( .A(instr[7]), .B(n1856), .D(n1857), .C(n1828), .Y(n1855) );
  INVX1 U2324 ( .A(ramwe), .Y(n2131) );
  AO222X1 U2325 ( .A(dph_current[6]), .B(n616), .C(dptr_inc[14]), .D(n99), .E(
        n1307), .F(temp[6]), .Y(n1623) );
  AO44X1 U2326 ( .A(n903), .B(n1876), .C(instr[7]), .D(n446), .E(n1945), .F(
        instr[4]), .G(n736), .H(n1948), .Y(n751) );
  OAI31XL U2327 ( .A(n1689), .B(n2068), .C(n63), .D(n2086), .Y(n1876) );
  INVX1 U2328 ( .A(n1123), .Y(n2086) );
  NAND21X1 U2329 ( .B(instr[5]), .A(instr[4]), .Y(n793) );
  NAND21X1 U2330 ( .B(n121), .A(n446), .Y(n1026) );
  OR3XL U2331 ( .A(n121), .B(n809), .C(n1117), .Y(n506) );
  OAI22X1 U2332 ( .A(n1695), .B(n124), .C(n431), .D(n716), .Y(n954) );
  NOR4XL U2333 ( .A(n1696), .B(n1697), .C(n908), .D(n1674), .Y(n1695) );
  NOR3XL U2334 ( .A(n2030), .B(instr[3]), .C(n1692), .Y(n1697) );
  OAI222XL U2335 ( .A(n2042), .B(n1159), .C(n1698), .D(n2099), .E(n1699), .F(
        n2037), .Y(n1696) );
  AOI21BBXL U2336 ( .B(n1864), .C(n1865), .A(n104), .Y(n890) );
  XNOR2XL U2337 ( .A(n2105), .B(n1958), .Y(n1864) );
  XNOR2XL U2338 ( .A(n442), .B(n2188), .Y(n1865) );
  OAI22X1 U2339 ( .A(n124), .B(n953), .C(n431), .D(n952), .Y(n1296) );
  AND4X1 U2340 ( .A(n1668), .B(n1669), .C(n1667), .D(n2034), .Y(n952) );
  AOI211X1 U2341 ( .C(n1892), .D(n2189), .A(n951), .B(n2018), .Y(n953) );
  NOR2X1 U2342 ( .A(n908), .B(n1674), .Y(n1668) );
  OAI211X1 U2343 ( .C(n1627), .D(n1628), .A(n69), .B(n933), .Y(n1618) );
  NOR4XL U2344 ( .A(instr[2]), .B(instr[0]), .C(n1911), .D(n16), .Y(n1627) );
  AOI21X1 U2345 ( .B(n1629), .C(n1630), .A(n445), .Y(n1628) );
  AOI32X1 U2346 ( .A(instr[6]), .B(n960), .C(n2193), .D(n1631), .E(n1116), .Y(
        n1630) );
  OAI211X1 U2347 ( .C(n902), .D(n1061), .A(n1062), .B(phase[0]), .Y(n615) );
  OA22X1 U2348 ( .A(n1868), .B(n1869), .C(n63), .D(n1870), .Y(n887) );
  AOI32X1 U2349 ( .A(n1124), .B(n63), .C(instr[1]), .D(n1682), .E(n1957), .Y(
        n1869) );
  GEN2XL U2350 ( .D(n2039), .E(n1871), .C(n2188), .B(n1957), .A(n1872), .Y(
        n1870) );
  AOI222XL U2351 ( .A(n445), .B(n57), .C(n2188), .D(n1873), .E(n1948), .F(
        n2106), .Y(n1868) );
  AO22X1 U2352 ( .A(n1424), .B(pc_o[8]), .C(pc_i[8]), .D(n1905), .Y(n639) );
  AO21X1 U2353 ( .B(n923), .C(phase[1]), .A(n1571), .Y(n643) );
  NOR2X1 U2354 ( .A(n2085), .B(n2188), .Y(n902) );
  INVX1 U2355 ( .A(ramdatao[7]), .Y(n2130) );
  INVX1 U2356 ( .A(ramdatao[5]), .Y(n2141) );
  NOR2X1 U2357 ( .A(n2095), .B(instr[6]), .Y(n1123) );
  NOR3XL U2358 ( .A(n2039), .B(instr[3]), .C(n2095), .Y(n1822) );
  NAND4X1 U2359 ( .A(phase[0]), .B(n1124), .C(n1753), .D(n442), .Y(n1662) );
  OAI211X1 U2360 ( .C(n2194), .D(n1699), .A(n1754), .B(n1755), .Y(n1753) );
  OAI21X1 U2361 ( .B(n1631), .C(n1682), .A(n2194), .Y(n1754) );
  NAND2X1 U2362 ( .A(dec_cop[6]), .B(n116), .Y(n1212) );
  INVX1 U2363 ( .A(ramdatao[6]), .Y(n2136) );
  ENOX1 U2364 ( .A(n2053), .B(n88), .C(N11852), .D(n1309), .Y(dph_current[0])
         );
  MUX2X1 U2365 ( .D0(n254), .D1(n253), .S(n119), .Y(N11852) );
  MUX4X1 U2366 ( .D0(dph_reg[0]), .D1(dph_reg[8]), .D2(dph_reg[16]), .D3(
        dph_reg[24]), .S0(n436), .S1(n434), .Y(n254) );
  MUX4X1 U2367 ( .D0(dph_reg[32]), .D1(dph_reg[40]), .D2(dph_reg[48]), .D3(
        dph_reg[56]), .S0(n436), .S1(n434), .Y(n253) );
  AND2X1 U2368 ( .A(dec_cop[7]), .B(n115), .Y(n1213) );
  NAND2X1 U2369 ( .A(dec_cop[4]), .B(n116), .Y(n1214) );
  AOI22X1 U2370 ( .A(n10), .B(n1116), .C(n2193), .D(n1839), .Y(n1115) );
  OAI222XL U2371 ( .A(n1159), .B(n2098), .C(n1681), .D(n2082), .E(n737), .F(
        n2093), .Y(n1676) );
  AOI22X1 U2372 ( .A(n2194), .B(n1124), .C(n1331), .D(n121), .Y(n1681) );
  INVX1 U2373 ( .A(temp2_comb[0]), .Y(n1225) );
  AOI221XL U2374 ( .A(n9), .B(n901), .C(n449), .D(n2193), .E(n1123), .Y(n1692)
         );
  AOI22X1 U2375 ( .A(n1955), .B(n2190), .C(n15), .D(instr[4]), .Y(n1699) );
  NAND2X1 U2376 ( .A(dec_cop[3]), .B(n115), .Y(n1228) );
  AOI211X1 U2377 ( .C(n1594), .D(n1489), .A(n1670), .B(n1671), .Y(n1669) );
  NOR4XL U2378 ( .A(n446), .B(instr[3]), .C(n1672), .D(n16), .Y(n1671) );
  AOI21X1 U2379 ( .B(n2193), .C(instr[1]), .A(n1673), .Y(n1672) );
  OAI21BBX1 U2380 ( .A(n1687), .B(n1946), .C(n1685), .Y(n951) );
  OAI21X1 U2381 ( .B(n2042), .C(n1689), .A(n89), .Y(n1687) );
  AOI221XL U2382 ( .A(n1594), .B(instr[3]), .C(n1686), .D(n891), .E(n1670), 
        .Y(n1685) );
  AOI32X1 U2383 ( .A(instr[6]), .B(n442), .C(n1911), .D(n1167), .E(n2085), .Y(
        n1698) );
  INVX1 U2384 ( .A(n922), .Y(n715) );
  AOI211X1 U2385 ( .C(n1676), .D(n369), .A(n1677), .B(n1678), .Y(n1675) );
  OAI31XL U2386 ( .A(n916), .B(instr[6]), .C(n2190), .D(n1679), .Y(n1678) );
  NAND2X1 U2387 ( .A(n1116), .B(instr[1]), .Y(n896) );
  GEN2XL U2388 ( .D(n1945), .E(n1895), .C(n743), .B(n433), .A(n813), .Y(n834)
         );
  OAI31XL U2389 ( .A(n929), .B(n737), .C(n2084), .D(n930), .Y(n813) );
  NAND3X1 U2390 ( .A(n64), .B(n89), .C(n931), .Y(n929) );
  OAI22X1 U2391 ( .A(n2068), .B(n1954), .C(n431), .D(n736), .Y(n931) );
  AO222X1 U2392 ( .A(dph_current[7]), .B(n616), .C(dptr_inc[15]), .D(n99), .E(
        n1307), .F(temp[7]), .Y(n1632) );
  ENOX1 U2393 ( .A(n2130), .B(n88), .C(N11845), .D(n1309), .Y(dph_current[7])
         );
  MUX2X1 U2394 ( .D0(n268), .D1(n267), .S(n118), .Y(N11845) );
  MUX2X1 U2395 ( .D0(ramsfraddr[6]), .D1(n1454), .S(waitstaten), .Y(
        ramsfraddr_comb[6]) );
  MUX2X1 U2396 ( .D0(ramsfraddr[5]), .D1(n1711), .S(n2184), .Y(
        ramsfraddr_comb[5]) );
  AND2X1 U2397 ( .A(dec_cop[2]), .B(n116), .Y(n1207) );
  INVX1 U2398 ( .A(acc[4]), .Y(n2140) );
  AND2X1 U2399 ( .A(dec_cop[5]), .B(n115), .Y(n1209) );
  ENOX1 U2400 ( .A(n2120), .B(n88), .C(N11850), .D(n1309), .Y(dph_current[2])
         );
  MUX2X1 U2401 ( .D0(n258), .D1(n257), .S(n119), .Y(N11850) );
  MUX4X1 U2402 ( .D0(dph_reg[2]), .D1(dph_reg[10]), .D2(dph_reg[18]), .D3(
        dph_reg[26]), .S0(N346), .S1(N347), .Y(n258) );
  MUX4X1 U2403 ( .D0(dph_reg[34]), .D1(dph_reg[42]), .D2(dph_reg[50]), .D3(
        dph_reg[58]), .S0(N346), .S1(N347), .Y(n257) );
  ENOX1 U2404 ( .A(n2064), .B(n88), .C(N11851), .D(n1309), .Y(dph_current[1])
         );
  MUX2X1 U2405 ( .D0(n256), .D1(n255), .S(n118), .Y(N11851) );
  MUX4X1 U2406 ( .D0(dph_reg[1]), .D1(dph_reg[9]), .D2(dph_reg[17]), .D3(
        dph_reg[25]), .S0(N346), .S1(n434), .Y(n256) );
  MUX4X1 U2407 ( .D0(dph_reg[33]), .D1(dph_reg[41]), .D2(dph_reg[49]), .D3(
        dph_reg[57]), .S0(N346), .S1(n434), .Y(n255) );
  MUX2X1 U2408 ( .D0(ramsfraddr[7]), .D1(n1455), .S(n450), .Y(
        ramsfraddr_comb[7]) );
  AOI21X1 U2409 ( .B(n1956), .C(instr[6]), .A(n1683), .Y(n1849) );
  INVX1 U2410 ( .A(temp2_comb[7]), .Y(n2160) );
  AOI33X1 U2411 ( .A(n1852), .B(n1958), .C(n1331), .D(n1167), .E(n1956), .F(
        n10), .Y(n1851) );
  OAI21X1 U2412 ( .B(instr[6]), .C(n449), .A(n2082), .Y(n1852) );
  NOR2X1 U2413 ( .A(n2092), .B(instr[3]), .Y(n1636) );
  NAND3X1 U2414 ( .A(n1636), .B(interrupt), .C(n1688), .Y(n1667) );
  NOR3XL U2415 ( .A(n445), .B(instr[1]), .C(n2097), .Y(n1688) );
  AOI21X1 U2416 ( .B(n2188), .C(instr[4]), .A(n1124), .Y(n1872) );
  INVX1 U2417 ( .A(temp[4]), .Y(n2155) );
  INVX1 U2418 ( .A(temp[3]), .Y(n2152) );
  NAND2X1 U2419 ( .A(dec_cop[1]), .B(n115), .Y(n1206) );
  INVX1 U2420 ( .A(n778), .Y(n794) );
  OAI31XL U2421 ( .A(instr[7]), .B(n2100), .C(n2033), .D(n2081), .Y(n778) );
  NAND32X1 U2422 ( .B(n121), .C(n2088), .A(n1947), .Y(n1757) );
  MUX2X1 U2423 ( .D0(n1423), .D1(n21), .S(pc_o[1]), .Y(n740) );
  NAND21X1 U2424 ( .B(n1456), .A(temp2_comb[0]), .Y(n640) );
  INVX1 U2425 ( .A(acc[6]), .Y(n1556) );
  INVX1 U2426 ( .A(acc[0]), .Y(n783) );
  ENOX1 U2427 ( .A(n2128), .B(n88), .C(N11849), .D(n1309), .Y(dph_current[3])
         );
  MUX2X1 U2428 ( .D0(n260), .D1(n259), .S(n118), .Y(N11849) );
  MUX4X1 U2429 ( .D0(dph_reg[3]), .D1(dph_reg[11]), .D2(dph_reg[19]), .D3(
        dph_reg[27]), .S0(N346), .S1(N347), .Y(n260) );
  MUX4X1 U2430 ( .D0(dph_reg[35]), .D1(dph_reg[43]), .D2(dph_reg[51]), .D3(
        dph_reg[59]), .S0(N346), .S1(N347), .Y(n259) );
  OAI22X1 U2431 ( .A(instr[7]), .B(n2033), .C(n917), .D(n2030), .Y(n913) );
  INVX1 U2432 ( .A(dec_accop[10]), .Y(n2116) );
  INVX1 U2433 ( .A(temp[2]), .Y(n1964) );
  INVX1 U2434 ( .A(temp[6]), .Y(n1965) );
  INVX1 U2435 ( .A(temp[1]), .Y(n2151) );
  INVX1 U2436 ( .A(temp[0]), .Y(n2129) );
  INVX1 U2437 ( .A(temp[5]), .Y(n2157) );
  AOI221XL U2438 ( .A(n2023), .B(memaddr[9]), .C(memdatai[1]), .D(n1136), .E(
        n1148), .Y(n1147) );
  OAI22X1 U2439 ( .A(n1913), .B(n1138), .C(n2022), .D(n2173), .Y(n1148) );
  NAND21X1 U2440 ( .B(N343), .A(n1959), .Y(n786) );
  NAND21X1 U2441 ( .B(N344), .A(N343), .Y(n784) );
  NAND21X1 U2442 ( .B(N343), .A(N344), .Y(n1562) );
  NAND21X1 U2443 ( .B(n1959), .A(N343), .Y(n1606) );
  AO2222XL U2444 ( .A(multemp2[7]), .B(n501), .C(b[5]), .D(n504), .E(n408), 
        .F(n1949), .G(n503), .H(n493), .Y(N12482) );
  AO2222XL U2445 ( .A(b[3]), .B(n504), .C(n503), .D(n494), .E(n414), .F(n1949), 
        .G(multemp2[5]), .H(n501), .Y(N12480) );
  AO2222XL U2446 ( .A(b[1]), .B(n504), .C(n503), .D(n495), .E(n421), .F(n1949), 
        .G(multemp2[3]), .H(n501), .Y(N12478) );
  AO2222XL U2447 ( .A(b[6]), .B(n504), .C(n503), .D(n496), .E(n405), .F(n1949), 
        .G(multemp2[8]), .H(n501), .Y(N12483) );
  AO2222XL U2448 ( .A(b[4]), .B(n504), .C(n503), .D(n497), .E(n411), .F(n1949), 
        .G(multemp2[6]), .H(n501), .Y(N12481) );
  AO2222XL U2449 ( .A(b[2]), .B(n504), .C(n503), .D(n498), .E(n417), .F(n1949), 
        .G(multemp2[4]), .H(n501), .Y(N12479) );
  AO2222XL U2450 ( .A(b[0]), .B(n504), .C(n503), .D(n502), .E(n425), .F(n1949), 
        .G(multemp2[2]), .H(n501), .Y(N12477) );
  MUX2X1 U2451 ( .D0(n788), .D1(n787), .S(N345), .Y(n789) );
  OA2222XL U2452 ( .A(n783), .B(n786), .C(n2127), .D(n784), .E(n1967), .F(
        n1562), .G(n2154), .H(n1606), .Y(n788) );
  OA2222XL U2453 ( .A(n786), .B(n2140), .C(n784), .D(n2159), .E(n1562), .F(
        n1556), .G(n1966), .H(n1606), .Y(n787) );
  INVX1 U2454 ( .A(n835), .Y(n849) );
  NAND43X1 U2455 ( .B(p2sel), .C(n1898), .D(n843), .A(n1897), .Y(n835) );
  ENOX1 U2456 ( .A(n2134), .B(n88), .C(N11848), .D(n1309), .Y(dph_current[4])
         );
  MUX2X1 U2457 ( .D0(n262), .D1(n261), .S(n119), .Y(N11848) );
  MUX4X1 U2458 ( .D0(dph_reg[4]), .D1(dph_reg[12]), .D2(dph_reg[20]), .D3(
        dph_reg[28]), .S0(N346), .S1(N347), .Y(n262) );
  MUX4X1 U2459 ( .D0(dph_reg[36]), .D1(dph_reg[44]), .D2(dph_reg[52]), .D3(
        dph_reg[60]), .S0(N346), .S1(N347), .Y(n261) );
  ENOX1 U2460 ( .A(n2141), .B(n88), .C(N11847), .D(n1309), .Y(dph_current[5])
         );
  MUX2X1 U2461 ( .D0(n264), .D1(n263), .S(n118), .Y(N11847) );
  MUX4X1 U2462 ( .D0(dph_reg[5]), .D1(dph_reg[13]), .D2(dph_reg[21]), .D3(
        dph_reg[29]), .S0(N346), .S1(N347), .Y(n264) );
  MUX4X1 U2463 ( .D0(dph_reg[37]), .D1(dph_reg[45]), .D2(dph_reg[53]), .D3(
        dph_reg[61]), .S0(n436), .S1(N347), .Y(n263) );
  INVX1 U2464 ( .A(N344), .Y(n1959) );
  BUFX3 U2465 ( .A(pc_o[5]), .Y(memaddr[5]) );
  OAI22XL U2466 ( .A(n1130), .B(n1547), .C(n1135), .D(n461), .Y(N12720) );
  AOI221XL U2467 ( .A(n2023), .B(pc_o[14]), .C(memdatai[6]), .D(n1136), .E(
        n1137), .Y(n1135) );
  OAI22X1 U2468 ( .A(n1900), .B(n1138), .C(n2022), .D(n2168), .Y(n1137) );
  OAI22XL U2469 ( .A(n1130), .B(n1544), .C(n1139), .D(n461), .Y(N12719) );
  AOI221XL U2470 ( .A(n2023), .B(n49), .C(memdatai[5]), .D(n1136), .E(n1140), 
        .Y(n1139) );
  OAI22X1 U2471 ( .A(n1901), .B(n1138), .C(n2022), .D(n2169), .Y(n1140) );
  OAI22XL U2472 ( .A(n1130), .B(n1541), .C(n1141), .D(n460), .Y(N12718) );
  AOI221XL U2473 ( .A(n2023), .B(pc_o[12]), .C(memdatai[4]), .D(n1136), .E(
        n1142), .Y(n1141) );
  OAI22X1 U2474 ( .A(n1902), .B(n1138), .C(n2022), .D(n2170), .Y(n1142) );
  OAI22XL U2475 ( .A(n1130), .B(n1534), .C(n1143), .D(n460), .Y(N12717) );
  AOI221XL U2476 ( .A(n2023), .B(memaddr[11]), .C(memdatai[3]), .D(n1136), .E(
        n1144), .Y(n1143) );
  OAI22X1 U2477 ( .A(n1903), .B(n1138), .C(n2022), .D(n2171), .Y(n1144) );
  OAI22XL U2478 ( .A(n1130), .B(n1343), .C(n1145), .D(n461), .Y(N12716) );
  AOI221XL U2479 ( .A(n2023), .B(pc_o[10]), .C(memdatai[2]), .D(n1136), .E(
        n1146), .Y(n1145) );
  OAI22X1 U2480 ( .A(n1912), .B(n1138), .C(n2022), .D(n2172), .Y(n1146) );
  INVX1 U2481 ( .A(n489), .Y(n501) );
  NAND32X1 U2482 ( .B(n2113), .C(n491), .A(n1926), .Y(n489) );
  ENOX1 U2483 ( .A(n2136), .B(n88), .C(N11846), .D(n1309), .Y(dph_current[6])
         );
  MUX2X1 U2484 ( .D0(n266), .D1(n265), .S(n119), .Y(N11846) );
  MUX4X1 U2485 ( .D0(dph_reg[6]), .D1(dph_reg[14]), .D2(dph_reg[22]), .D3(
        dph_reg[30]), .S0(n285), .S1(n287), .Y(n266) );
  MUX4X1 U2486 ( .D0(dph_reg[38]), .D1(dph_reg[46]), .D2(dph_reg[54]), .D3(
        dph_reg[62]), .S0(n285), .S1(n287), .Y(n265) );
  INVX1 U2487 ( .A(n492), .Y(n503) );
  NAND32X1 U2488 ( .B(n2112), .C(n491), .A(n1925), .Y(n492) );
  NAND3X1 U2489 ( .A(ramsfraddr[3]), .B(ramsfraddr[4]), .C(n1007), .Y(n1013)
         );
  OAI221X1 U2490 ( .A(n2144), .B(n1342), .C(n795), .D(n2001), .E(n456), .Y(
        N12491) );
  INVX1 U2491 ( .A(p2[6]), .Y(n2144) );
  OAI221X1 U2492 ( .A(n2143), .B(n1342), .C(n795), .D(n2000), .E(n456), .Y(
        N12492) );
  INVX1 U2493 ( .A(p2[7]), .Y(n2143) );
  OAI221X1 U2494 ( .A(n2146), .B(n1342), .C(n795), .D(n2003), .E(n456), .Y(
        N12489) );
  INVX1 U2495 ( .A(p2[4]), .Y(n2146) );
  OAI221X1 U2496 ( .A(n2147), .B(n1342), .C(n2004), .D(n795), .E(n456), .Y(
        N12488) );
  INVX1 U2497 ( .A(p2[3]), .Y(n2147) );
  OAI221X1 U2498 ( .A(n2145), .B(n1342), .C(n2002), .D(n795), .E(n456), .Y(
        N12490) );
  INVX1 U2499 ( .A(p2[5]), .Y(n2145) );
  INVX1 U2500 ( .A(phase[3]), .Y(n1954) );
  OAI22X1 U2501 ( .A(n1168), .B(n2001), .C(n1170), .D(n1190), .Y(N12706) );
  EORX1 U2502 ( .A(n1191), .B(ac), .C(n1192), .D(n1179), .Y(n1190) );
  NAND21X1 U2503 ( .B(n1927), .A(n1187), .Y(n1191) );
  AOI32X1 U2504 ( .A(n2116), .B(n2115), .C(N11555), .D(dec_accop[10]), .E(
        n2063), .Y(n1192) );
  OAI22X1 U2505 ( .A(n1168), .B(n2005), .C(n1169), .D(n1170), .Y(N12711) );
  AOI211X1 U2506 ( .C(ov), .D(n1171), .A(n1172), .B(n1173), .Y(n1169) );
  NAND3X1 U2507 ( .A(n1185), .B(n1186), .C(n1187), .Y(n1171) );
  AOI21X1 U2508 ( .B(n1174), .C(n1175), .A(n1176), .Y(n1173) );
  ENOX1 U2509 ( .A(n685), .B(n2005), .C(gf0), .D(n685), .Y(n1881) );
  AND2X1 U2510 ( .A(n686), .B(n452), .Y(n685) );
  ENOX1 U2511 ( .A(n687), .B(n2006), .C(f1), .D(n687), .Y(n1883) );
  ENOX1 U2512 ( .A(n688), .B(n2004), .C(n688), .D(dps[3]), .Y(n1884) );
  NOR2X1 U2513 ( .A(n459), .B(n2074), .Y(n688) );
  ENOX1 U2514 ( .A(n687), .B(n2002), .C(f0), .D(n687), .Y(n1882) );
  MUX4X1 U2515 ( .D0(dph_reg[7]), .D1(dph_reg[15]), .D2(dph_reg[23]), .D3(
        dph_reg[31]), .S0(n285), .S1(n287), .Y(n268) );
  MUX4X1 U2516 ( .D0(dph_reg[39]), .D1(dph_reg[47]), .D2(dph_reg[55]), .D3(
        dph_reg[63]), .S0(n285), .S1(n287), .Y(n267) );
  NAND21X1 U2517 ( .B(state[0]), .A(n680), .Y(n1078) );
  AND2X1 U2518 ( .A(phase0_ff), .B(n451), .Y(newinstr) );
  NOR21XL U2519 ( .B(phase[4]), .A(n723), .Y(N684) );
  NOR21XL U2520 ( .B(n394), .A(n1345), .Y(N12484) );
  AOI22X1 U2521 ( .A(n1346), .B(n1347), .C(n1949), .D(ramdatao[7]), .Y(n1345)
         );
  OAI21BBX1 U2522 ( .A(n1348), .B(b[7]), .C(n1349), .Y(n1346) );
  AOI33X1 U2523 ( .A(finishdiv), .B(n1925), .C(n1607), .D(multemp2[9]), .E(
        finishmul), .F(n1926), .Y(n1349) );
  NOR2X1 U2524 ( .A(state[1]), .B(state[2]), .Y(n680) );
  NOR32XL U2525 ( .B(n389), .C(n102), .A(newinstrlock), .Y(N689) );
  AND2X1 U2526 ( .A(state[1]), .B(n393), .Y(N589) );
  AND2X1 U2527 ( .A(state[2]), .B(n393), .Y(N590) );
  AOI21BX1 U2528 ( .C(n830), .B(n829), .A(n398), .Y(N12730) );
  AOI221XL U2529 ( .A(n2024), .B(pc_o[7]), .C(n1071), .D(ramdatai[7]), .E(
        n1067), .Y(n829) );
  OAI221X1 U2530 ( .A(n1566), .B(n2090), .C(n828), .D(n1087), .E(n1063), .Y(
        n830) );
  OAI222XL U2531 ( .A(n2161), .B(n1068), .C(n2160), .D(n2027), .E(n2054), .F(
        n1069), .Y(n1067) );
  AOI21BX1 U2532 ( .C(n857), .B(n856), .A(n397), .Y(N12728) );
  AOI221XL U2533 ( .A(n2024), .B(n2186), .C(n1071), .D(ramdatai[5]), .E(n1080), 
        .Y(n856) );
  OAI221X1 U2534 ( .A(n847), .B(n2090), .C(n1901), .D(n1087), .E(n1077), .Y(
        n857) );
  OAI222XL U2535 ( .A(n2157), .B(n1068), .C(n2158), .D(n2027), .E(n2056), .F(
        n1069), .Y(n1080) );
  AOI21BX1 U2536 ( .C(n864), .B(n863), .A(n399), .Y(N12727) );
  AOI221XL U2537 ( .A(n2024), .B(memaddr[4]), .C(n1071), .D(ramdatai[4]), .E(
        n1084), .Y(n863) );
  OAI221X1 U2538 ( .A(n853), .B(n2090), .C(n1902), .D(n1087), .E(n1081), .Y(
        n864) );
  OAI222XL U2539 ( .A(n2155), .B(n1068), .C(n2156), .D(n2027), .E(n2057), .F(
        n1069), .Y(n1084) );
  AOI21BX1 U2540 ( .C(n875), .B(n874), .A(n399), .Y(N12726) );
  AOI221XL U2541 ( .A(n2024), .B(pc_o[3]), .C(n1071), .D(ramdatai[3]), .E(
        n1088), .Y(n874) );
  OAI221X1 U2542 ( .A(n1533), .B(n2090), .C(n1903), .D(n1087), .E(n1085), .Y(
        n875) );
  OAI222XL U2543 ( .A(n2152), .B(n1068), .C(n2153), .D(n2027), .E(n2058), .F(
        n1069), .Y(n1088) );
  AOI21BX1 U2544 ( .C(n939), .B(n938), .A(n399), .Y(N12729) );
  AOI221XL U2545 ( .A(n2024), .B(pc_o[6]), .C(n1071), .D(ramdatai[6]), .E(
        n1076), .Y(n938) );
  OAI221X1 U2546 ( .A(n841), .B(n2090), .C(n1900), .D(n1087), .E(n1073), .Y(
        n939) );
  OAI222XL U2547 ( .A(n1965), .B(n1068), .C(n2139), .D(n2027), .E(n2055), .F(
        n1069), .Y(n1076) );
  AOI21BX1 U2548 ( .C(n1101), .B(n1099), .A(n399), .Y(N12723) );
  OAI221X1 U2549 ( .A(n1131), .B(n2090), .C(n1091), .D(n1087), .E(n1100), .Y(
        n1101) );
  AOI221XL U2550 ( .A(n2024), .B(N1761), .C(pc_i[8]), .D(n1095), .E(n1102), 
        .Y(n1099) );
  AOI221XL U2551 ( .A(n2026), .B(temp[0]), .C(n1089), .D(temp2_comb[0]), .E(
        n21), .Y(n1100) );
  AOI31X1 U2552 ( .A(n1090), .B(n1092), .C(n566), .D(n397), .Y(N12725) );
  AOI221XL U2553 ( .A(n1089), .B(temp2_comb[2]), .C(n2026), .D(temp[2]), .E(
        n1093), .Y(n1092) );
  OA22X1 U2554 ( .A(n1912), .B(n1087), .C(n865), .D(n2090), .Y(n566) );
  AOI22X1 U2555 ( .A(n1071), .B(ramdatai[2]), .C(n1072), .D(memdatai[2]), .Y(
        n1090) );
  AOI31X1 U2556 ( .A(n1096), .B(n1097), .C(n985), .D(n399), .Y(N12724) );
  OA22X1 U2557 ( .A(n43), .B(n1094), .C(n1069), .D(n984), .Y(n985) );
  AOI221XL U2558 ( .A(n2026), .B(temp[1]), .C(n1089), .D(temp2_comb[1]), .E(
        n22), .Y(n1096) );
  AOI221XL U2559 ( .A(n1071), .B(ramdatai[1]), .C(n1072), .D(memdatai[1]), .E(
        n1098), .Y(n1097) );
  INVX1 U2560 ( .A(phase[4]), .Y(n767) );
  AOI31X1 U2561 ( .A(n745), .B(n1940), .C(n747), .D(n684), .Y(n744) );
  AOI22X1 U2562 ( .A(phase[2]), .B(n750), .C(phase[3]), .D(n751), .Y(n745) );
  AOI221XL U2563 ( .A(n432), .B(n748), .C(n102), .D(n749), .E(codefetch_s), 
        .Y(n747) );
  NOR2X1 U2564 ( .A(n1023), .B(n1024), .Y(N12976) );
  AOI21X1 U2565 ( .B(waitcnt[0]), .C(waitcnt[1]), .A(waitcnt[2]), .Y(n1023) );
  NOR2X1 U2566 ( .A(n1025), .B(n1024), .Y(N12975) );
  XNOR2XL U2567 ( .A(waitcnt[1]), .B(waitcnt[0]), .Y(n1025) );
  NOR2X1 U2568 ( .A(waitcnt[0]), .B(n1024), .Y(N12974) );
  INVX1 U2569 ( .A(idle_r), .Y(n1953) );
  INVX1 U2570 ( .A(temp[7]), .Y(n2161) );
  AOI22X1 U2571 ( .A(n1072), .B(memdatai[7]), .C(intvect[4]), .D(n22), .Y(
        n1063) );
  AOI22X1 U2572 ( .A(n1072), .B(memdatai[5]), .C(intvect[2]), .D(n22), .Y(
        n1077) );
  AOI22X1 U2573 ( .A(n1072), .B(memdatai[4]), .C(intvect[1]), .D(n21), .Y(
        n1081) );
  AOI22X1 U2574 ( .A(n1072), .B(memdatai[3]), .C(intvect[0]), .D(n21), .Y(
        n1085) );
  AOI22X1 U2575 ( .A(n1072), .B(memdatai[6]), .C(intvect[3]), .D(n21), .Y(
        n1073) );
  AND3X1 U2576 ( .A(n653), .B(acc[3]), .C(n2014), .Y(n1522) );
  OAI21X1 U2577 ( .B(idle_r), .C(stop_r), .A(n695), .Y(n693) );
  INVX1 U2578 ( .A(n499), .Y(n502) );
  MUX2AXL U2579 ( .D0(N13345), .D1(n1556), .S(N13353), .Y(n499) );
  NAND5XL U2580 ( .A(n1944), .B(n1962), .C(n832), .D(n831), .E(ramsfraddr[5]), 
        .Y(n795) );
  INVX1 U2581 ( .A(n1000), .Y(n832) );
  OAI31XL U2582 ( .A(n1177), .B(n1178), .C(n1179), .D(n1180), .Y(n1172) );
  NAND42X1 U2583 ( .C(b[3]), .D(b[4]), .A(n1181), .B(n1182), .Y(n1180) );
  XNOR2XL U2584 ( .A(n1184), .B(n2062), .Y(n1177) );
  NOR3XL U2585 ( .A(b[5]), .B(b[7]), .C(b[6]), .Y(n1181) );
  INVX1 U2586 ( .A(p2[0]), .Y(n2150) );
  INVX1 U2587 ( .A(p2[1]), .Y(n2149) );
  AOI21BX1 U2588 ( .C(cpu_hold), .B(d_hold), .A(cpu_resume_fff), .Y(n726) );
  INVX1 U2589 ( .A(p2[2]), .Y(n2148) );
  AO21X1 U2590 ( .B(N343), .C(N344), .A(n1908), .Y(n196) );
  INVX1 U2591 ( .A(n1305), .Y(n1974) );
  OAI221X1 U2592 ( .A(n2054), .B(n78), .C(n1267), .D(n17), .E(n1306), .Y(n1305) );
  AOI222XL U2593 ( .A(N11793), .B(n1269), .C(N11827), .D(n1270), .E(N11810), 
        .F(n1271), .Y(n1306) );
  OA21X1 U2594 ( .B(N343), .C(n1959), .A(n2036), .Y(n197) );
  INVX1 U2595 ( .A(n1312), .Y(n1976) );
  OAI221X1 U2596 ( .A(n2056), .B(n78), .C(n65), .D(n47), .E(n1313), .Y(n1312)
         );
  AOI222XL U2597 ( .A(N11791), .B(n87), .C(N11825), .D(n98), .E(N11808), .F(
        n111), .Y(n1313) );
  INVX1 U2598 ( .A(n1310), .Y(n1975) );
  OAI221X1 U2599 ( .A(n2055), .B(n78), .C(n65), .D(n41), .E(n1311), .Y(n1310)
         );
  AOI222XL U2600 ( .A(N11792), .B(n87), .C(N11826), .D(n1270), .E(N11809), .F(
        n1271), .Y(n1311) );
  OAI211X1 U2601 ( .C(n1154), .D(n431), .A(n1155), .B(n1107), .Y(n1136) );
  OAI31XL U2602 ( .A(n886), .B(n1156), .C(n919), .D(n102), .Y(n1155) );
  NOR42XL U2603 ( .C(n1158), .D(n716), .A(n1162), .B(n1163), .Y(n1154) );
  OAI21X1 U2604 ( .B(ramsfraddr[7]), .C(n1153), .A(n658), .Y(n1132) );
  NAND2X1 U2605 ( .A(state[0]), .B(n680), .Y(n684) );
  INVX1 U2606 ( .A(n1288), .Y(n2032) );
  OAI221X1 U2607 ( .A(memaddr[0]), .B(n78), .C(n65), .D(n37), .E(n1289), .Y(
        n1288) );
  AOI222XL U2608 ( .A(N1761), .B(n87), .C(memaddr[0]), .D(n98), .E(n37), .F(
        n111), .Y(n1289) );
  INVX1 U2609 ( .A(n1278), .Y(n1984) );
  OAI221X1 U2610 ( .A(n2061), .B(n78), .C(n65), .D(n23), .E(n1279), .Y(n1278)
         );
  AOI222XL U2611 ( .A(N11783), .B(n87), .C(N11817), .D(n1270), .E(N11800), .F(
        n1271), .Y(n1279) );
  INVX1 U2612 ( .A(n1318), .Y(n1979) );
  OAI221X1 U2613 ( .A(n2059), .B(n78), .C(n65), .D(n27), .E(n1319), .Y(n1318)
         );
  AOI222XL U2614 ( .A(N11788), .B(n87), .C(N11822), .D(n98), .E(N11805), .F(
        n111), .Y(n1319) );
  INVX1 U2615 ( .A(n1316), .Y(n1978) );
  OAI221X1 U2616 ( .A(n2058), .B(n78), .C(n65), .D(n29), .E(n1317), .Y(n1316)
         );
  AOI222XL U2617 ( .A(N11789), .B(n87), .C(N11823), .D(n1270), .E(N11806), .F(
        n1271), .Y(n1317) );
  INVX1 U2618 ( .A(n1314), .Y(n1977) );
  OAI221X1 U2619 ( .A(n2057), .B(n78), .C(n65), .D(n35), .E(n1315), .Y(n1314)
         );
  AOI222XL U2620 ( .A(N11790), .B(n87), .C(N11824), .D(n98), .E(N11807), .F(
        n111), .Y(n1315) );
  INVX1 U2621 ( .A(N345), .Y(n2118) );
  INVX1 U2622 ( .A(stop_r), .Y(n1960) );
  OAI21X1 U2623 ( .B(n1110), .C(n1111), .A(n102), .Y(n1104) );
  GEN2XL U2624 ( .D(n1116), .E(n1117), .C(n1118), .B(n1119), .A(n1120), .Y(
        n1110) );
  OAI222XL U2625 ( .A(n89), .B(n1112), .C(n1113), .D(n1114), .E(n2190), .F(
        n1115), .Y(n1111) );
  OAI31XL U2626 ( .A(n2039), .B(n16), .C(n1121), .D(n1122), .Y(n1120) );
  AOI211X1 U2627 ( .C(instr[2]), .D(n2039), .A(instr[3]), .B(n901), .Y(n1113)
         );
  INVX1 U2628 ( .A(state[0]), .Y(n1059) );
  NAND31X1 U2629 ( .C(n1153), .A(ramsfraddr[7]), .B(n452), .Y(n1130) );
  AOI21X1 U2630 ( .B(n102), .C(n743), .A(n1897), .Y(n1109) );
  NAND2X1 U2631 ( .A(n1898), .B(instr[4]), .Y(n1069) );
  NAND2X1 U2632 ( .A(n433), .B(n1164), .Y(n1151) );
  OAI21X1 U2633 ( .B(n1165), .C(n2093), .A(n1166), .Y(n1164) );
  AOI22X1 U2634 ( .A(n1167), .B(n120), .C(n1948), .D(n2190), .Y(n1165) );
  NOR4XL U2635 ( .A(b[2]), .B(b[1]), .C(b[0]), .D(n1183), .Y(n1182) );
  AOI21X1 U2636 ( .B(n121), .C(n1124), .A(n2190), .Y(n1121) );
  INVX1 U2637 ( .A(pdmode), .Y(n2009) );
  AND2X1 U2638 ( .A(n1152), .B(n102), .Y(n1128) );
  OAI21BX1 U2639 ( .C(n972), .B(n1789), .A(n432), .Y(n1819) );
  NAND3X1 U2640 ( .A(n1012), .B(n1923), .C(ramsfraddr[5]), .Y(n1347) );
  OAI21X1 U2641 ( .B(n1788), .C(n1605), .A(n102), .Y(n1820) );
  INVX1 U2642 ( .A(finishdiv), .Y(n2112) );
  INVX1 U2643 ( .A(finishmul), .Y(n2113) );
  AND2X1 U2644 ( .A(cpu_resume_ff1), .B(n457), .Y(N13380) );
  NOR2X1 U2645 ( .A(n2115), .B(dec_accop[10]), .Y(n1178) );
  OAI22AX1 U2646 ( .D(ckcon[7]), .C(n1029), .A(n2130), .B(n1030), .Y(N12972)
         );
  NOR2X1 U2647 ( .A(phase[2]), .B(n432), .Y(n1817) );
  NAND3X1 U2648 ( .A(n2071), .B(n2119), .C(ramsfraddr[2]), .Y(n1003) );
  NAND3X1 U2649 ( .A(ramsfraddr[0]), .B(n2119), .C(ramsfraddr[2]), .Y(n1004)
         );
  INVXL U2650 ( .A(n1419), .Y(n1432) );
  MUX2X2 U2651 ( .D0(pc_o[4]), .D1(n1481), .S(n146), .Y(memaddr_comb[4]) );
  MUX2X1 U2652 ( .D0(memaddr[0]), .D1(n1476), .S(n146), .Y(memaddr_comb[0]) );
  AND3XL U2653 ( .A(n1840), .B(n1272), .C(n1248), .Y(n1273) );
  NAND43X1 U2654 ( .B(n1272), .C(n1078), .D(interrupt), .A(n2009), .Y(n1079)
         );
  OA21XL U2655 ( .B(n1272), .C(n1075), .A(n680), .Y(n1074) );
  NAND21XL U2656 ( .B(n1272), .A(n1052), .Y(n1058) );
  NAND21XL U2657 ( .B(pdmode), .A(n1272), .Y(n1050) );
  NAND21X2 U2658 ( .B(n766), .A(n765), .Y(n1272) );
  MUX2X2 U2659 ( .D0(pc_o[2]), .D1(n1478), .S(n146), .Y(memaddr_comb[2]) );
  NAND21XL U2660 ( .B(n2118), .A(n1402), .Y(n1604) );
  NAND21X2 U2661 ( .B(N345), .A(n1402), .Y(n1304) );
  NAND32X2 U2662 ( .B(n692), .C(n579), .A(n691), .Y(n1402) );
  INVX1 U2663 ( .A(n1404), .Y(n1413) );
  AND2XL U2664 ( .A(n389), .B(n1300), .Y(N11498) );
  NAND42XL U2665 ( .C(n472), .D(n469), .A(n466), .B(n465), .Y(n382) );
  INVX1 U2666 ( .A(n382), .Y(n451) );
  INVX1 U2667 ( .A(n382), .Y(n450) );
  AOI22XL U2668 ( .A(sfrdatai[7]), .B(n1915), .C(n1391), .D(n970), .Y(n1385)
         );
  INVX2 U2669 ( .A(sfrdatai[7]), .Y(n1564) );
  MUX2XL U2670 ( .D0(pc_o[9]), .D1(n1500), .S(n145), .Y(memaddr_comb[9]) );
  MUX2XL U2671 ( .D0(pc_o[10]), .D1(n1501), .S(n145), .Y(memaddr_comb[10]) );
  MUX2XL U2672 ( .D0(pc_o[8]), .D1(n1491), .S(n145), .Y(memaddr_comb[8]) );
  MUX2XL U2673 ( .D0(pc_o[7]), .D1(n1485), .S(n145), .Y(memaddr_comb[7]) );
  MUX2X1 U2674 ( .D0(pc_o[3]), .D1(n1479), .S(n145), .Y(memaddr_comb[3]) );
  MUX2X1 U2675 ( .D0(memaddr[5]), .D1(n1483), .S(n145), .Y(memaddr_comb[5]) );
  MUX2XL U2676 ( .D0(memaddr[1]), .D1(n1477), .S(n146), .Y(memaddr_comb[1]) );
  AND2X1 U2677 ( .A(sfrwe_r), .B(n2184), .Y(sfrwe) );
  NAND21X2 U2678 ( .B(n786), .A(n1530), .Y(n694) );
  NAND31X2 U2679 ( .C(n698), .A(n697), .B(n694), .Y(n699) );
  NOR21X2 U2680 ( .B(n702), .A(n701), .Y(n703) );
  NAND32X1 U2681 ( .B(n762), .C(n761), .A(n760), .Y(n764) );
  OA2222X1 U2682 ( .A(n1913), .B(n1539), .C(n1456), .D(n2126), .E(n759), .F(
        n1553), .G(n1537), .H(n758), .Y(n760) );
  AOI221X1 U2683 ( .A(n754), .B(n172), .C(n1530), .D(n1433), .E(n753), .Y(n759) );
  OAI22XL U2684 ( .A(n1294), .B(n1293), .C(n1292), .D(n1773), .Y(n1295) );
  INVXL U2685 ( .A(n1300), .Y(n1294) );
  AOI211XL U2686 ( .C(n1530), .D(n1529), .A(n1528), .B(n1527), .Y(n1538) );
  OAI22XL U2687 ( .A(n1130), .B(n1352), .C(n1147), .D(n460), .Y(N12715) );
  OAI211XL U2688 ( .C(n1352), .D(n1510), .A(n540), .B(n539), .Y(n983) );
  INVX2 U2689 ( .A(sfrdatai[1]), .Y(n1352) );
  NOR21XL U2690 ( .B(n1301), .A(n1293), .Y(n995) );
  MUX2X2 U2691 ( .D0(n764), .D1(n983), .S(n1904), .Y(n1301) );
  NAND21XL U2692 ( .B(n398), .A(n1475), .Y(n804) );
  NAND21XL U2693 ( .B(n1475), .A(n388), .Y(n805) );
  NAND21XL U2694 ( .B(n1475), .A(n976), .Y(n958) );
  NAND21X2 U2695 ( .B(n690), .A(n689), .Y(n691) );
  MUX2IX2 U2696 ( .D0(n682), .D1(n679), .S(N345), .Y(n689) );
  AO2222X1 U2697 ( .A(n1529), .B(n1519), .C(n677), .D(n1302), .E(n1433), .F(
        n741), .G(n1415), .H(n669), .Y(n682) );
  AO2222X1 U2698 ( .A(n1529), .B(n1574), .C(n677), .D(n1554), .E(n1433), .F(
        n1419), .G(n1415), .H(n1404), .Y(n679) );
  OAI22XL U2699 ( .A(n1322), .B(n1308), .C(n1562), .D(n1304), .Y(n1390) );
  AOI22XL U2700 ( .A(sfrdatai[4]), .B(n1915), .C(n967), .D(n1391), .Y(n1465)
         );
  AO2222XL U2701 ( .A(ramdatao[7]), .B(n148), .C(n961), .D(n959), .E(n958), 
        .F(pc_o[15]), .G(p2[7]), .H(n149), .Y(n1506) );
  AO2222XL U2702 ( .A(n148), .B(ramdatao[6]), .C(n850), .D(n959), .E(n958), 
        .F(memaddr[14]), .G(p2[6]), .H(n149), .Y(n1505) );
  AO2222XL U2703 ( .A(n148), .B(ramdatao[5]), .C(n858), .D(n959), .E(n958), 
        .F(n49), .G(p2[5]), .H(n149), .Y(n1504) );
  AO2222XL U2704 ( .A(n148), .B(ramdatao[4]), .C(n867), .D(n959), .E(n958), 
        .F(memaddr[12]), .G(p2[4]), .H(n149), .Y(n1503) );
  AO2222XL U2705 ( .A(n148), .B(ramdatao[3]), .C(n876), .D(n959), .E(n958), 
        .F(memaddr[11]), .G(p2[3]), .H(n149), .Y(n1502) );
  MAJ3X1 U2706 ( .A(N11541), .B(N11549), .C(N11522), .Y(n530) );
  MAJ3X1 U2707 ( .A(N11523), .B(N11542), .C(n530), .Y(
        add_1_root_add_5140_2_carry[2]) );
  NOR32X4 U2708 ( .B(n641), .C(n640), .A(n639), .Y(n704) );
  NOR21X4 U2709 ( .B(n700), .A(n699), .Y(n701) );
  NOR43X4 U2710 ( .B(n706), .C(n705), .D(n704), .A(n703), .Y(n709) );
  INVX8 U2711 ( .A(n1086), .Y(n708) );
  MUX2IX4 U2712 ( .D0(n709), .D1(n708), .S(n1904), .Y(n1300) );
  MUX2IX4 U2713 ( .D0(idle), .D1(n1300), .S(n981), .Y(n738) );
  MUX2IX4 U2714 ( .D0(stop), .D1(n1301), .S(n981), .Y(n765) );
  MAJ3X1 U2715 ( .A(n1568), .B(n1354), .C(n1353), .Y(n1535) );
  MAJ3X1 U2716 ( .A(n1568), .B(n1535), .C(n161), .Y(n1542) );
  MAJ3X1 U2717 ( .A(n1568), .B(n1542), .C(n162), .Y(n1545) );
  MAJ3X1 U2718 ( .A(n1568), .B(n1545), .C(n163), .Y(n1548) );
  MAJ3X1 U2719 ( .A(n1568), .B(n1548), .C(n164), .Y(n1567) );
  MAJ3X1 U2720 ( .A(n1568), .B(n1567), .C(n165), .Y(n1570) );
  XNOR2XL U2721 ( .A(pc_o[15]), .B(add_5280_3_carry_15_), .Y(N11810) );
  OR2X1 U2722 ( .A(add_5280_3_carry_14_), .B(memaddr[14]), .Y(
        add_5280_3_carry_15_) );
  XNOR2XL U2723 ( .A(add_5280_3_carry_14_), .B(pc_o[14]), .Y(N11809) );
  OR2X1 U2724 ( .A(add_5280_3_carry_13_), .B(n49), .Y(add_5280_3_carry_14_) );
  XNOR2XL U2725 ( .A(add_5280_3_carry_13_), .B(n49), .Y(N11808) );
  OR2X1 U2726 ( .A(add_5280_3_carry_12_), .B(memaddr[12]), .Y(
        add_5280_3_carry_13_) );
  XNOR2XL U2727 ( .A(add_5280_3_carry_12_), .B(memaddr[12]), .Y(N11807) );
  OR2X1 U2728 ( .A(add_5280_3_carry_11_), .B(memaddr[11]), .Y(
        add_5280_3_carry_12_) );
  XNOR2XL U2729 ( .A(add_5280_3_carry_11_), .B(memaddr[11]), .Y(N11806) );
  OR2X1 U2730 ( .A(add_5280_3_carry_10_), .B(pc_o[10]), .Y(
        add_5280_3_carry_11_) );
  XNOR2XL U2731 ( .A(add_5280_3_carry_10_), .B(pc_o[10]), .Y(N11805) );
  OR2X1 U2732 ( .A(add_5280_3_carry_9_), .B(memaddr[9]), .Y(
        add_5280_3_carry_10_) );
  XNOR2XL U2733 ( .A(add_5280_3_carry_9_), .B(memaddr[9]), .Y(N11804) );
  OR2X1 U2734 ( .A(add_5280_3_carry_8_), .B(pc_o[8]), .Y(add_5280_3_carry_9_)
         );
  XNOR2XL U2735 ( .A(add_5280_3_carry_8_), .B(memaddr[8]), .Y(N11803) );
  OR2X1 U2736 ( .A(add_5280_3_carry_7_), .B(pc_o[7]), .Y(add_5280_3_carry_8_)
         );
  XNOR2XL U2737 ( .A(add_5280_3_carry_7_), .B(n2185), .Y(N11802) );
  OR2X1 U2738 ( .A(add_5280_3_carry_6_), .B(pc_o[6]), .Y(add_5280_3_carry_7_)
         );
  XNOR2XL U2739 ( .A(add_5280_3_carry_6_), .B(pc_o[6]), .Y(N11801) );
  OR2X1 U2740 ( .A(add_5280_3_carry_5_), .B(pc_o[5]), .Y(add_5280_3_carry_6_)
         );
  XNOR2XL U2741 ( .A(add_5280_3_carry_5_), .B(pc_o[5]), .Y(N11800) );
  OR2X1 U2742 ( .A(add_5280_3_carry_4_), .B(memaddr[4]), .Y(
        add_5280_3_carry_5_) );
  XNOR2XL U2743 ( .A(add_5280_3_carry_4_), .B(memaddr[4]), .Y(N11799) );
  OR2X1 U2744 ( .A(add_5280_3_carry_3_), .B(memaddr[3]), .Y(
        add_5280_3_carry_4_) );
  XNOR2XL U2745 ( .A(add_5280_3_carry_3_), .B(pc_o[3]), .Y(N11798) );
  OR2X1 U2746 ( .A(add_5280_3_carry_2_), .B(memaddr[2]), .Y(
        add_5280_3_carry_3_) );
  XNOR2XL U2747 ( .A(add_5280_3_carry_2_), .B(pc_o[2]), .Y(N11797) );
  OR2X1 U2748 ( .A(N1761), .B(pc_o[1]), .Y(add_5280_3_carry_2_) );
  XNOR2XL U2749 ( .A(pc_o[0]), .B(memaddr[1]), .Y(N11796) );
  XNOR2XL U2750 ( .A(pc_o[15]), .B(add_5280_4_carry[15]), .Y(N11827) );
  OR2X1 U2751 ( .A(add_5280_4_carry[14]), .B(pc_o[14]), .Y(
        add_5280_4_carry[15]) );
  XNOR2XL U2752 ( .A(add_5280_4_carry[14]), .B(memaddr[14]), .Y(N11826) );
  OR2X1 U2753 ( .A(add_5280_4_carry[13]), .B(n49), .Y(add_5280_4_carry[14]) );
  XNOR2XL U2754 ( .A(add_5280_4_carry[13]), .B(n49), .Y(N11825) );
  OR2X1 U2755 ( .A(add_5280_4_carry[12]), .B(pc_o[12]), .Y(
        add_5280_4_carry[13]) );
  XNOR2XL U2756 ( .A(add_5280_4_carry[12]), .B(pc_o[12]), .Y(N11824) );
  OR2X1 U2757 ( .A(add_5280_4_carry[11]), .B(pc_o[11]), .Y(
        add_5280_4_carry[12]) );
  XNOR2XL U2758 ( .A(add_5280_4_carry[11]), .B(pc_o[11]), .Y(N11823) );
  OR2X1 U2759 ( .A(add_5280_4_carry[10]), .B(memaddr[10]), .Y(
        add_5280_4_carry[11]) );
  XNOR2XL U2760 ( .A(add_5280_4_carry[10]), .B(memaddr[10]), .Y(N11822) );
  OR2X1 U2761 ( .A(add_5280_4_carry[9]), .B(pc_o[9]), .Y(add_5280_4_carry[10])
         );
  XNOR2XL U2762 ( .A(add_5280_4_carry[9]), .B(pc_o[9]), .Y(N11821) );
  OR2X1 U2763 ( .A(add_5280_4_carry[8]), .B(pc_o[8]), .Y(add_5280_4_carry[9])
         );
  XNOR2XL U2764 ( .A(add_5280_4_carry[8]), .B(pc_o[8]), .Y(N11820) );
  OR2X1 U2765 ( .A(add_5280_4_carry[7]), .B(pc_o[7]), .Y(add_5280_4_carry[8])
         );
  XNOR2XL U2766 ( .A(add_5280_4_carry[7]), .B(n2185), .Y(N11819) );
  OR2X1 U2767 ( .A(add_5280_4_carry[6]), .B(pc_o[6]), .Y(add_5280_4_carry[7])
         );
  XNOR2XL U2768 ( .A(add_5280_4_carry[6]), .B(memaddr[6]), .Y(N11818) );
  OR2X1 U2769 ( .A(add_5280_4_carry[5]), .B(memaddr[5]), .Y(
        add_5280_4_carry[6]) );
  XNOR2XL U2770 ( .A(add_5280_4_carry[5]), .B(n2186), .Y(N11817) );
  OR2X1 U2771 ( .A(add_5280_4_carry[4]), .B(pc_o[4]), .Y(add_5280_4_carry[5])
         );
  XNOR2XL U2772 ( .A(add_5280_4_carry[4]), .B(pc_o[4]), .Y(N11816) );
  OR2X1 U2773 ( .A(add_5280_4_carry[3]), .B(pc_o[3]), .Y(add_5280_4_carry[4])
         );
  XNOR2XL U2774 ( .A(add_5280_4_carry[3]), .B(memaddr[3]), .Y(N11815) );
  OR2X1 U2775 ( .A(pc_o[1]), .B(pc_o[2]), .Y(add_5280_4_carry[3]) );
  XNOR2XL U2776 ( .A(pc_o[1]), .B(memaddr[2]), .Y(N11814) );
  XOR2X1 U2777 ( .A(pc_o[15]), .B(add_5280_2_carry[15]), .Y(N11793) );
  AND2X1 U2778 ( .A(pc_o[14]), .B(add_5280_2_carry[14]), .Y(
        add_5280_2_carry[15]) );
  XOR2X1 U2779 ( .A(add_5280_2_carry[14]), .B(pc_o[14]), .Y(N11792) );
  AND2X1 U2780 ( .A(pc_o[13]), .B(add_5280_2_carry[13]), .Y(
        add_5280_2_carry[14]) );
  XOR2X1 U2781 ( .A(add_5280_2_carry[13]), .B(pc_o[13]), .Y(N11791) );
  AND2X1 U2782 ( .A(pc_o[12]), .B(add_5280_2_carry[12]), .Y(
        add_5280_2_carry[13]) );
  XOR2X1 U2783 ( .A(add_5280_2_carry[12]), .B(pc_o[12]), .Y(N11790) );
  AND2X1 U2784 ( .A(pc_o[11]), .B(add_5280_2_carry[11]), .Y(
        add_5280_2_carry[12]) );
  XOR2X1 U2785 ( .A(add_5280_2_carry[11]), .B(pc_o[11]), .Y(N11789) );
  AND2X1 U2786 ( .A(pc_o[10]), .B(add_5280_2_carry[10]), .Y(
        add_5280_2_carry[11]) );
  XOR2X1 U2787 ( .A(add_5280_2_carry[10]), .B(pc_o[10]), .Y(N11788) );
  AND2X1 U2788 ( .A(pc_o[9]), .B(add_5280_2_carry[9]), .Y(add_5280_2_carry[10]) );
  XOR2X1 U2789 ( .A(add_5280_2_carry[9]), .B(pc_o[9]), .Y(N11787) );
  AND2X1 U2790 ( .A(pc_o[8]), .B(add_5280_2_carry[8]), .Y(add_5280_2_carry[9])
         );
  XOR2X1 U2791 ( .A(add_5280_2_carry[8]), .B(pc_o[8]), .Y(N11786) );
  AND2X1 U2792 ( .A(pc_o[7]), .B(add_5280_2_carry[7]), .Y(add_5280_2_carry[8])
         );
  XOR2X1 U2793 ( .A(add_5280_2_carry[7]), .B(pc_o[7]), .Y(N11785) );
  AND2X1 U2794 ( .A(pc_o[6]), .B(add_5280_2_carry[6]), .Y(add_5280_2_carry[7])
         );
  XOR2X1 U2795 ( .A(add_5280_2_carry[6]), .B(pc_o[6]), .Y(N11784) );
  AND2X1 U2796 ( .A(pc_o[5]), .B(add_5280_2_carry[5]), .Y(add_5280_2_carry[6])
         );
  XOR2X1 U2797 ( .A(add_5280_2_carry[5]), .B(pc_o[5]), .Y(N11783) );
  AND2X1 U2798 ( .A(pc_o[4]), .B(add_5280_2_carry[4]), .Y(add_5280_2_carry[5])
         );
  XOR2X1 U2799 ( .A(add_5280_2_carry[4]), .B(pc_o[4]), .Y(N11782) );
  AND2X1 U2800 ( .A(memaddr[3]), .B(add_5280_2_carry[3]), .Y(
        add_5280_2_carry[4]) );
  XOR2X1 U2801 ( .A(add_5280_2_carry[3]), .B(pc_o[3]), .Y(N11781) );
  AND2X1 U2802 ( .A(memaddr[2]), .B(pc_o[1]), .Y(add_5280_2_carry[3]) );
  XOR2X1 U2803 ( .A(pc_o[1]), .B(pc_o[2]), .Y(N11780) );
  XOR2X1 U2804 ( .A(n2185), .B(add_1469_carry[7]), .Y(N1768) );
  AND2X1 U2805 ( .A(pc_o[6]), .B(add_1469_carry[6]), .Y(add_1469_carry[7]) );
  XOR2X1 U2806 ( .A(add_1469_carry[6]), .B(memaddr[6]), .Y(N1767) );
  AND2X1 U2807 ( .A(pc_o[5]), .B(add_1469_carry[5]), .Y(add_1469_carry[6]) );
  XOR2X1 U2808 ( .A(add_1469_carry[5]), .B(memaddr[5]), .Y(N1766) );
  AND2X1 U2809 ( .A(memaddr[4]), .B(add_1469_carry[4]), .Y(add_1469_carry[5])
         );
  XOR2X1 U2810 ( .A(add_1469_carry[4]), .B(pc_o[4]), .Y(N1765) );
  AND2X1 U2811 ( .A(pc_o[3]), .B(add_1469_carry[3]), .Y(add_1469_carry[4]) );
  XOR2X1 U2812 ( .A(add_1469_carry[3]), .B(pc_o[3]), .Y(N1764) );
  AND2X1 U2813 ( .A(pc_o[2]), .B(memaddr[1]), .Y(add_1469_carry[3]) );
  XOR2X1 U2814 ( .A(pc_o[1]), .B(pc_o[2]), .Y(N1763) );
  XNOR2XL U2815 ( .A(N12776), .B(add_5526_carry_7_), .Y(N12817) );
  OR2X1 U2816 ( .A(add_5526_carry_6_), .B(N12775), .Y(add_5526_carry_7_) );
  XNOR2XL U2817 ( .A(add_5526_carry_6_), .B(N12775), .Y(N12816) );
  OR2X1 U2818 ( .A(add_5526_carry_5_), .B(N12774), .Y(add_5526_carry_6_) );
  XNOR2XL U2819 ( .A(add_5526_carry_5_), .B(N12774), .Y(N12815) );
  OR2X1 U2820 ( .A(add_5526_carry_4_), .B(N12773), .Y(add_5526_carry_5_) );
  XNOR2XL U2821 ( .A(add_5526_carry_4_), .B(N12773), .Y(N12814) );
  OR2X1 U2822 ( .A(add_5526_carry_3_), .B(N12772), .Y(add_5526_carry_4_) );
  XNOR2XL U2823 ( .A(add_5526_carry_3_), .B(N12772), .Y(N12813) );
  OR2X1 U2824 ( .A(add_5526_carry_2_), .B(N12771), .Y(add_5526_carry_3_) );
  XNOR2XL U2825 ( .A(add_5526_carry_2_), .B(N12771), .Y(N12812) );
  OR2X1 U2826 ( .A(N12769), .B(N12770), .Y(add_5526_carry_2_) );
  XNOR2XL U2827 ( .A(N12769), .B(N12770), .Y(N12811) );
  AND2X1 U2828 ( .A(b[0]), .B(acc[0]), .Y(N14336) );
  AND2X1 U2829 ( .A(b[1]), .B(acc[0]), .Y(N14337) );
  AND2X1 U2830 ( .A(b[2]), .B(n112), .Y(N14338) );
  AND2X1 U2831 ( .A(b[3]), .B(n112), .Y(N14339) );
  AND2X1 U2832 ( .A(b[4]), .B(n112), .Y(N14340) );
  AND2X1 U2833 ( .A(b[5]), .B(n112), .Y(N14341) );
  AND2X1 U2834 ( .A(b[6]), .B(n112), .Y(N14342) );
  AND2X1 U2835 ( .A(n112), .B(b[7]), .Y(N14343) );
  AND2X1 U2836 ( .A(b[0]), .B(acc[1]), .Y(N14344) );
  AND2X1 U2837 ( .A(b[1]), .B(acc[1]), .Y(N14345) );
  AND2X1 U2838 ( .A(b[2]), .B(acc[1]), .Y(N14346) );
  AND2X1 U2839 ( .A(b[3]), .B(acc[1]), .Y(N14347) );
  AND2X1 U2840 ( .A(b[4]), .B(n106), .Y(N14348) );
  AND2X1 U2841 ( .A(b[5]), .B(n106), .Y(N14349) );
  AND2X1 U2842 ( .A(b[6]), .B(n106), .Y(N14350) );
  AND2X1 U2843 ( .A(n106), .B(b[7]), .Y(N14351) );
  INVX1 U2844 ( .A(N12769), .Y(N12810) );
  MAJ3X1 U2848 ( .A(N11545), .B(N11526), .C(N11555), .Y(n2180) );
endmodule


module mcu51_cpu_a0_DW01_add_7 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;

  wire   [7:1] carry;

  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(SUM[8]), .SO(SUM[7]) );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  XOR2X1 U1 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
  AND2X1 U2 ( .A(A[0]), .B(B[0]), .Y(carry[1]) );
endmodule


module mcu51_cpu_a0_DW01_add_8 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;

  wire   [7:1] carry;

  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(SUM[8]), .SO(SUM[7]) );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  AND2X1 U1 ( .A(A[0]), .B(B[0]), .Y(carry[1]) );
  XOR2X1 U2 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
endmodule


module mcu51_cpu_a0_DW01_inc_2 ( A, SUM );
  input [15:0] A;
  output [15:0] SUM;

  wire   [15:2] carry;

  HAD1X1 U1_1_14 ( .A(A[14]), .B(carry[14]), .CO(carry[15]), .SO(SUM[14]) );
  HAD1X1 U1_1_13 ( .A(A[13]), .B(carry[13]), .CO(carry[14]), .SO(SUM[13]) );
  HAD1X1 U1_1_12 ( .A(A[12]), .B(carry[12]), .CO(carry[13]), .SO(SUM[12]) );
  HAD1X1 U1_1_11 ( .A(A[11]), .B(carry[11]), .CO(carry[12]), .SO(SUM[11]) );
  HAD1X1 U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .SO(SUM[10]) );
  HAD1X1 U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .SO(SUM[9]) );
  HAD1X1 U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .SO(SUM[8]) );
  HAD1X1 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .SO(SUM[7]) );
  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  XOR2X1 U1 ( .A(carry[15]), .B(A[15]), .Y(SUM[15]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module mcu51_cpu_a0_DW01_inc_1 ( A, SUM );
  input [15:0] A;
  output [15:0] SUM;

  wire   [15:2] carry;

  HAD1X1 U1_1_14 ( .A(A[14]), .B(carry[14]), .CO(carry[15]), .SO(SUM[14]) );
  HAD1X1 U1_1_13 ( .A(A[13]), .B(carry[13]), .CO(carry[14]), .SO(SUM[13]) );
  HAD1X1 U1_1_12 ( .A(A[12]), .B(carry[12]), .CO(carry[13]), .SO(SUM[12]) );
  HAD1X1 U1_1_11 ( .A(A[11]), .B(carry[11]), .CO(carry[12]), .SO(SUM[11]) );
  HAD1X1 U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .SO(SUM[10]) );
  HAD1X1 U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .SO(SUM[9]) );
  HAD1X1 U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .SO(SUM[8]) );
  HAD1X1 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .SO(SUM[7]) );
  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  XOR2X1 U1 ( .A(carry[15]), .B(A[15]), .Y(SUM[15]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module mcu51_cpu_a0_DW01_inc_0 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  HAD1X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .SO(SUM[6]) );
  HAD1X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .SO(SUM[5]) );
  HAD1X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .SO(SUM[4]) );
  HAD1X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .SO(SUM[3]) );
  HAD1X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .SO(SUM[2]) );
  HAD1X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .SO(SUM[1]) );
  XOR2X1 U1 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module mcu51_cpu_a0_DW01_sub_1 ( A, B, CI, DIFF, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9;
  wire   [7:1] carry;

  FAD1X1 U2_6 ( .A(A[6]), .B(n5), .CI(carry[6]), .CO(carry[7]), .SO(DIFF[6])
         );
  FAD1X1 U2_5 ( .A(A[5]), .B(n8), .CI(carry[5]), .CO(carry[6]), .SO(DIFF[5])
         );
  FAD1X1 U2_4 ( .A(A[4]), .B(n4), .CI(carry[4]), .CO(carry[5]), .SO(DIFF[4])
         );
  FAD1X1 U2_3 ( .A(A[3]), .B(n7), .CI(carry[3]), .CO(carry[4]), .SO(DIFF[3])
         );
  FAD1X1 U2_2 ( .A(A[2]), .B(n3), .CI(carry[2]), .CO(carry[3]), .SO(DIFF[2])
         );
  FAD1X1 U2_1 ( .A(A[1]), .B(n6), .CI(carry[1]), .CO(carry[2]), .SO(DIFF[1])
         );
  INVX1 U1 ( .A(B[2]), .Y(n3) );
  INVX1 U2 ( .A(B[3]), .Y(n7) );
  INVX1 U3 ( .A(B[4]), .Y(n4) );
  INVX1 U4 ( .A(B[5]), .Y(n8) );
  INVX1 U5 ( .A(B[1]), .Y(n6) );
  NAND21X1 U6 ( .B(n2), .A(n1), .Y(carry[1]) );
  INVX1 U7 ( .A(A[0]), .Y(n1) );
  INVX1 U8 ( .A(B[6]), .Y(n5) );
  INVX1 U9 ( .A(B[0]), .Y(n2) );
  XOR2X1 U10 ( .A(B[0]), .B(A[0]), .Y(DIFF[0]) );
  AOI21X1 U11 ( .B(carry[7]), .C(A[7]), .A(n9), .Y(DIFF[8]) );
  AOI21BBXL U12 ( .B(A[7]), .C(carry[7]), .A(B[7]), .Y(n9) );
endmodule


module mcu51_cpu_a0_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9;
  wire   [8:1] carry;

  FAD1X1 U2_7 ( .A(A[7]), .B(n2), .CI(carry[7]), .CO(carry[8]), .SO(DIFF[7])
         );
  FAD1X1 U2_6 ( .A(A[6]), .B(n6), .CI(carry[6]), .CO(carry[7]), .SO(DIFF[6])
         );
  FAD1X1 U2_5 ( .A(A[5]), .B(n9), .CI(carry[5]), .CO(carry[6]), .SO(DIFF[5])
         );
  FAD1X1 U2_4 ( .A(A[4]), .B(n5), .CI(carry[4]), .CO(carry[5]), .SO(DIFF[4])
         );
  FAD1X1 U2_3 ( .A(A[3]), .B(n8), .CI(carry[3]), .CO(carry[4]), .SO(DIFF[3])
         );
  FAD1X1 U2_2 ( .A(A[2]), .B(n4), .CI(carry[2]), .CO(carry[3]), .SO(DIFF[2])
         );
  FAD1X1 U2_1 ( .A(A[1]), .B(n7), .CI(carry[1]), .CO(carry[2]), .SO(DIFF[1])
         );
  INVX1 U1 ( .A(B[2]), .Y(n4) );
  INVX1 U2 ( .A(B[3]), .Y(n8) );
  INVX1 U3 ( .A(B[4]), .Y(n5) );
  INVX1 U4 ( .A(B[5]), .Y(n9) );
  INVX1 U5 ( .A(B[6]), .Y(n6) );
  INVX1 U6 ( .A(B[1]), .Y(n7) );
  NAND21X1 U7 ( .B(n3), .A(n1), .Y(carry[1]) );
  INVX1 U8 ( .A(A[0]), .Y(n1) );
  INVX1 U9 ( .A(B[7]), .Y(n2) );
  INVX1 U10 ( .A(B[0]), .Y(n3) );
  XOR2X1 U11 ( .A(B[0]), .B(A[0]), .Y(DIFF[0]) );
  INVX1 U12 ( .A(carry[8]), .Y(DIFF[8]) );
endmodule


module mcu51_cpu_a0_DW01_add_0 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [15:1] carry;

  FAD1X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .SO(
        SUM[14]) );
  FAD1X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .SO(
        SUM[13]) );
  FAD1X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .SO(
        SUM[12]) );
  FAD1X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .SO(
        SUM[11]) );
  FAD1X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .SO(
        SUM[10]) );
  FAD1X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .SO(SUM[9])
         );
  FAD1X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .SO(SUM[8])
         );
  FAD1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .SO(SUM[7])
         );
  FAD1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .SO(SUM[6])
         );
  FAD1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .SO(SUM[5])
         );
  FAD1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .SO(SUM[4])
         );
  FAD1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .SO(SUM[3])
         );
  FAD1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .SO(SUM[2])
         );
  FAD1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .SO(SUM[1])
         );
  XOR3X1 U1_15 ( .A(A[15]), .B(B[15]), .C(carry[15]), .Y(SUM[15]) );
  XOR2X1 U1 ( .A(A[0]), .B(B[0]), .Y(SUM[0]) );
  INVX1 U2 ( .A(B[0]), .Y(n1) );
  NOR21XL U3 ( .B(A[0]), .A(n1), .Y(carry[1]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_3 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_4 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_5 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_6 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_7 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_8 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_9 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_10 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_11 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_12 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_13 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_14 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_15 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_16 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_17 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_18 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_19 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_20 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_21 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_22 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_23 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_24 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_25 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_26 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_27 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_28 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_29 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_30 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_31 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_32 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_33 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_34 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_35 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_36 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_37 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_38 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_39 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_40 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_41 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_42 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_43 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_44 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_45 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_46 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_47 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_48 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_49 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_50 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_51 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_52 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_53 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_54 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module SNPS_CLOCK_GATE_HIGH_mcu51_cpu_a0_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;


  CLKDLXL latch ( .CK(CLK), .E(EN), .SE(TE), .ECK(ENCLK) );
endmodule


module mpb_a0 ( i_rd, i_wr, wdat0, wdat1, addr0, addr1, r_i2c_attr, esfrm_oe, 
        esfrm_we, sfrack, esfrm_wdat, esfrm_adr, mcu_esfr_rdat, delay_rdat, 
        delay_rrdy, esfrm_rrdy, esfrm_rdat, channel_sel, r_pg0_sel, dma_w, 
        dma_r, dma_addr, dma_wdat, dma_ack, memaddr, memaddr_c, memwr, memrd, 
        memrd_c, cpurst, memdatao, memack, hit_xd, hit_xr, hit_ps, hit_ps_c, 
        idat_r, idat_w, idat_adr, idat_wdat, iram_ce, xram_ce, regx_re, 
        iram_we, xram_we, regx_we, iram_a, xram_a, iram_d, xram_d, iram_rdat, 
        xram_rdat, regx_rdat, bist_en, bist_wr, bist_adr, bist_wdat, bist_xram, 
        mclk, srstz );
  input [1:0] i_rd;
  input [1:0] i_wr;
  input [7:0] wdat0;
  input [7:0] wdat1;
  input [7:0] addr0;
  input [7:0] addr1;
  output [7:0] esfrm_wdat;
  output [6:0] esfrm_adr;
  input [7:0] mcu_esfr_rdat;
  input [7:0] delay_rdat;
  output [7:0] esfrm_rdat;
  input [3:0] r_pg0_sel;
  input [10:0] dma_addr;
  input [7:0] dma_wdat;
  input [15:0] memaddr;
  input [15:0] memaddr_c;
  input [7:0] memdatao;
  input [7:0] idat_adr;
  input [7:0] idat_wdat;
  output [10:0] iram_a;
  output [10:0] xram_a;
  output [7:0] iram_d;
  output [7:0] xram_d;
  input [7:0] iram_rdat;
  input [7:0] xram_rdat;
  input [7:0] regx_rdat;
  input [10:0] bist_adr;
  input [7:0] bist_wdat;
  input r_i2c_attr, delay_rrdy, channel_sel, dma_w, dma_r, memwr, memrd,
         memrd_c, cpurst, idat_r, idat_w, bist_en, bist_wr, bist_xram, mclk,
         srstz;
  output esfrm_oe, esfrm_we, sfrack, esfrm_rrdy, dma_ack, memack, hit_xd,
         hit_xr, hit_ps, hit_ps_c, iram_ce, xram_ce, regx_re, iram_we, xram_we,
         regx_we;
  wire   n229, dma_hit_x, pg0_rdwait, pg0_wrwait, N44, N45, r_pg0_rdrdy, N46,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228;
  wire   [1:0] xram_rdsel;

  DFFRQX1 r_pg0_rdrdy_reg ( .D(N46), .C(mclk), .XR(srstz), .Q(r_pg0_rdrdy) );
  DFFRQX1 xram_rdsel_reg_1_ ( .D(n191), .C(mclk), .XR(srstz), .Q(xram_rdsel[1]) );
  DFFRQX1 xram_rdsel_reg_0_ ( .D(n190), .C(mclk), .XR(srstz), .Q(xram_rdsel[0]) );
  DFFRQX1 pg0_rdwait_reg ( .D(N45), .C(mclk), .XR(srstz), .Q(pg0_rdwait) );
  DFFRQX1 pg0_wrwait_reg ( .D(N44), .C(mclk), .XR(srstz), .Q(pg0_wrwait) );
  BUFX3 U3 ( .A(n229), .Y(xram_a[1]) );
  NAND21X1 U4 ( .B(i_rd[1]), .A(n22), .Y(n21) );
  NAND21X1 U5 ( .B(n183), .A(n182), .Y(n188) );
  INVX1 U6 ( .A(n188), .Y(esfrm_oe) );
  INVX1 U7 ( .A(n29), .Y(n161) );
  NAND21X1 U8 ( .B(n131), .A(dma_addr[3]), .Y(n95) );
  NAND21X1 U9 ( .B(n131), .A(dma_addr[5]), .Y(n101) );
  NAND21X1 U10 ( .B(pg0_wrwait), .A(n23), .Y(n29) );
  NAND31X1 U11 ( .C(n184), .A(n186), .B(n185), .Y(n23) );
  INVX1 U12 ( .A(n139), .Y(n96) );
  OAI211X1 U13 ( .C(n52), .D(n66), .A(n72), .B(n51), .Y(xram_d[1]) );
  INVX1 U14 ( .A(n143), .Y(n102) );
  OAI2B11X1 U15 ( .D(dma_addr[1]), .C(n131), .A(n134), .B(n91), .Y(n229) );
  OAI2B11X1 U16 ( .D(dma_addr[4]), .C(n131), .A(n141), .B(n98), .Y(xram_a[4])
         );
  AND4X1 U17 ( .A(memaddr[11]), .B(memaddr[7]), .C(n211), .D(n212), .Y(hit_xr)
         );
  OA33X1 U18 ( .A(n161), .B(n167), .C(n160), .D(n159), .E(bist_en), .F(n158), 
        .Y(n3) );
  INVX1 U19 ( .A(n164), .Y(n4) );
  INVX1 U20 ( .A(n167), .Y(n5) );
  NAND2X1 U21 ( .A(r_pg0_sel[2]), .B(n19), .Y(n18) );
  INVX1 U22 ( .A(n18), .Y(n6) );
  INVX1 U23 ( .A(n18), .Y(n7) );
  INVX1 U24 ( .A(n20), .Y(n8) );
  OAI2B11X1 U25 ( .D(dma_addr[2]), .C(n131), .A(n137), .B(n92), .Y(xram_a[2])
         );
  BUFX3 U26 ( .A(bist_en), .Y(n192) );
  INVX1 U27 ( .A(n192), .Y(n9) );
  INVX1 U28 ( .A(n192), .Y(n10) );
  INVX1 U29 ( .A(n93), .Y(n11) );
  OA21X1 U30 ( .B(n140), .C(n126), .A(n11), .Y(n94) );
  INVXL U31 ( .A(n12), .Y(esfrm_adr[5]) );
  OAI2B11X1 U32 ( .D(dma_addr[6]), .C(n131), .A(n144), .B(n105), .Y(xram_a[6])
         );
  INVXL U33 ( .A(n155), .Y(n181) );
  NAND21XL U34 ( .B(n41), .A(n30), .Y(n156) );
  NAND21XL U35 ( .B(n161), .A(n30), .Y(n166) );
  AND2XL U36 ( .A(n181), .B(n41), .Y(n34) );
  AO22XL U37 ( .A(idat_adr[2]), .B(n136), .C(n149), .D(esfrm_adr[2]), .Y(n138)
         );
  AO22XL U38 ( .A(idat_adr[1]), .B(n136), .C(n149), .D(esfrm_adr[1]), .Y(n135)
         );
  OAI221XL U39 ( .A(n140), .B(n167), .C(n207), .D(n164), .E(n139), .Y(
        iram_a[3]) );
  AO21XL U40 ( .B(n177), .C(hit_xr), .A(n169), .Y(regx_we) );
  INVX1 U41 ( .A(n101), .Y(n13) );
  NAND43X1 U42 ( .B(n103), .C(n102), .D(n13), .A(n100), .Y(xram_a[5]) );
  NOR21XL U43 ( .B(memaddr[5]), .A(n128), .Y(n103) );
  INVX1 U44 ( .A(n95), .Y(n14) );
  NAND43X1 U45 ( .B(n97), .C(n96), .D(n14), .A(n94), .Y(xram_a[3]) );
  NOR21XL U46 ( .B(memaddr[3]), .A(n128), .Y(n97) );
  MUX2IXL U47 ( .D0(addr1[5]), .D1(addr0[5]), .S(n104), .Y(n12) );
  AO21XL U48 ( .B(n183), .C(n182), .A(pg0_rdwait), .Y(n39) );
  INVX1 U49 ( .A(n131), .Y(n112) );
  INVX1 U50 ( .A(i_wr[1]), .Y(n22) );
  INVX1 U51 ( .A(n166), .Y(n27) );
  INVX1 U52 ( .A(n126), .Y(n119) );
  INVX1 U53 ( .A(n164), .Y(n136) );
  INVX1 U54 ( .A(n167), .Y(n149) );
  NAND21X1 U55 ( .B(n162), .A(n88), .Y(n131) );
  AO21X1 U56 ( .B(n41), .C(n161), .A(n30), .Y(n155) );
  NAND21XL U57 ( .B(i_wr[0]), .A(n22), .Y(n185) );
  INVX4 U58 ( .A(n21), .Y(n104) );
  INVX1 U59 ( .A(n86), .Y(n88) );
  INVX1 U60 ( .A(n128), .Y(n111) );
  INVX1 U61 ( .A(n125), .Y(n118) );
  INVX1 U62 ( .A(n46), .Y(n64) );
  NAND32X1 U63 ( .B(bist_en), .C(n45), .A(n86), .Y(n46) );
  INVX1 U64 ( .A(n47), .Y(n45) );
  NAND21X1 U65 ( .B(bist_en), .A(n181), .Y(n126) );
  NAND21X1 U66 ( .B(bist_en), .A(n45), .Y(n66) );
  NAND21X1 U67 ( .B(bist_en), .A(n69), .Y(n167) );
  INVX1 U68 ( .A(n68), .Y(n69) );
  NAND21X1 U69 ( .B(bist_en), .A(n68), .Y(n164) );
  AO21X1 U70 ( .B(n69), .C(n43), .A(n171), .Y(N46) );
  AND2X1 U71 ( .A(n43), .B(n68), .Y(N45) );
  NAND21X1 U72 ( .B(n9), .A(bist_wdat[0]), .Y(n70) );
  NAND21X1 U73 ( .B(n10), .A(bist_wdat[1]), .Y(n72) );
  NAND21X1 U74 ( .B(n10), .A(bist_wdat[5]), .Y(n80) );
  NAND21X1 U75 ( .B(n9), .A(bist_wdat[4]), .Y(n78) );
  NAND21X1 U76 ( .B(n10), .A(bist_wdat[2]), .Y(n74) );
  NAND21X1 U77 ( .B(n10), .A(bist_wdat[3]), .Y(n76) );
  NAND21X1 U78 ( .B(n10), .A(bist_wr), .Y(n165) );
  INVX1 U79 ( .A(n195), .Y(n108) );
  INVX1 U80 ( .A(n48), .Y(n63) );
  NAND32X1 U81 ( .B(bist_en), .C(n86), .A(n47), .Y(n48) );
  INVX1 U82 ( .A(n90), .Y(esfrm_adr[0]) );
  INVXL U83 ( .A(n146), .Y(esfrm_adr[6]) );
  INVX1 U84 ( .A(n142), .Y(esfrm_adr[4]) );
  NOR21XL U85 ( .B(memaddr_c[3]), .A(n125), .Y(n93) );
  AOI21BBXL U86 ( .B(n12), .C(n126), .A(n99), .Y(n100) );
  NOR21XL U87 ( .B(memaddr_c[5]), .A(n125), .Y(n99) );
  INVX1 U88 ( .A(n39), .Y(n41) );
  OR2XL U89 ( .A(i_rd[0]), .B(i_rd[1]), .Y(n182) );
  INVX1 U90 ( .A(n159), .Y(n177) );
  NAND32X1 U91 ( .B(n88), .C(n162), .A(n87), .Y(n128) );
  AO21X1 U92 ( .B(n44), .C(n179), .A(n190), .Y(n86) );
  NAND21X1 U93 ( .B(n138), .A(n137), .Y(iram_a[2]) );
  OAI221XL U94 ( .A(n142), .B(n167), .C(n206), .D(n164), .E(n141), .Y(
        iram_a[4]) );
  NAND32X1 U95 ( .B(n162), .C(n87), .A(n86), .Y(n125) );
  NAND21X1 U96 ( .B(idat_r), .A(n163), .Y(n68) );
  INVX1 U97 ( .A(idat_w), .Y(n163) );
  OAI211X1 U98 ( .C(n191), .D(n3), .A(n175), .B(n174), .Y(xram_ce) );
  MUX3IX1 U99 ( .D0(n173), .D1(n172), .D2(bist_xram), .S0(n190), .S1(bist_en), 
        .Y(n174) );
  AND2X1 U100 ( .A(n191), .B(dma_hit_x), .Y(n173) );
  OAI31XL U101 ( .A(memaddr_c[15]), .B(memaddr_c[14]), .C(n193), .D(n191), .Y(
        n172) );
  INVX1 U102 ( .A(n31), .Y(n32) );
  OAI221XL U103 ( .A(n146), .B(n167), .C(n164), .D(n145), .E(n144), .Y(
        iram_a[6]) );
  INVX1 U104 ( .A(idat_adr[6]), .Y(n145) );
  OAI221X1 U105 ( .A(n12), .B(n167), .C(n205), .D(n164), .E(n143), .Y(
        iram_a[5]) );
  NAND32X1 U106 ( .B(n5), .C(bist_adr[8]), .A(n164), .Y(iram_a[8]) );
  OAI221X1 U107 ( .A(n197), .B(n126), .C(n198), .D(n10), .E(n117), .Y(
        xram_a[8]) );
  NAND21X1 U108 ( .B(n135), .A(n134), .Y(iram_a[1]) );
  OAI211X1 U109 ( .C(n153), .D(n164), .A(n167), .B(n152), .Y(iram_a[10]) );
  OAI211X1 U110 ( .C(n131), .D(n130), .A(n152), .B(n129), .Y(xram_a[10]) );
  NOR32XL U111 ( .B(n151), .C(n150), .A(n208), .Y(n153) );
  NAND21X1 U112 ( .B(n133), .A(n132), .Y(iram_a[0]) );
  AO22X1 U113 ( .A(idat_adr[0]), .B(n136), .C(n149), .D(esfrm_adr[0]), .Y(n133) );
  NAND21X1 U114 ( .B(n83), .A(n82), .Y(iram_d[6]) );
  AO22X1 U115 ( .A(idat_wdat[6]), .B(n136), .C(esfrm_wdat[6]), .D(n149), .Y(
        n83) );
  NAND21X1 U116 ( .B(n85), .A(n84), .Y(iram_d[7]) );
  AO22X1 U117 ( .A(idat_wdat[7]), .B(n136), .C(esfrm_wdat[7]), .D(n5), .Y(n85)
         );
  NAND21X1 U118 ( .B(n81), .A(n80), .Y(iram_d[5]) );
  AO22X1 U119 ( .A(idat_wdat[5]), .B(n136), .C(esfrm_wdat[5]), .D(n149), .Y(
        n81) );
  NAND21X1 U120 ( .B(n77), .A(n76), .Y(iram_d[3]) );
  AO22X1 U121 ( .A(idat_wdat[3]), .B(n4), .C(esfrm_wdat[3]), .D(n149), .Y(n77)
         );
  INVX1 U122 ( .A(n20), .Y(n30) );
  NAND21X1 U123 ( .B(n6), .A(n160), .Y(n20) );
  NAND21X1 U124 ( .B(n79), .A(n78), .Y(iram_d[4]) );
  AO22X1 U125 ( .A(idat_wdat[4]), .B(n136), .C(esfrm_wdat[4]), .D(n149), .Y(
        n79) );
  NAND21X1 U126 ( .B(n171), .A(n170), .Y(regx_re) );
  NAND43X1 U127 ( .B(n203), .C(n169), .D(n194), .A(n168), .Y(n170) );
  AND4X1 U128 ( .A(memaddr_c[9]), .B(memaddr_c[8]), .C(n190), .D(n191), .Y(
        n168) );
  INVX1 U129 ( .A(n127), .Y(n19) );
  NAND21X1 U130 ( .B(n75), .A(n74), .Y(iram_d[2]) );
  AO22X1 U131 ( .A(idat_wdat[2]), .B(n136), .C(esfrm_wdat[2]), .D(n149), .Y(
        n75) );
  NAND21X1 U132 ( .B(n71), .A(n70), .Y(iram_d[0]) );
  AO22X1 U133 ( .A(idat_wdat[0]), .B(n136), .C(n149), .D(esfrm_wdat[0]), .Y(
        n71) );
  NAND21X1 U134 ( .B(n73), .A(n72), .Y(iram_d[1]) );
  AO22X1 U135 ( .A(idat_wdat[1]), .B(n136), .C(esfrm_wdat[1]), .D(n149), .Y(
        n73) );
  INVX1 U136 ( .A(n157), .Y(n169) );
  NAND21XL U137 ( .B(n161), .A(n7), .Y(n157) );
  INVX1 U138 ( .A(n50), .Y(esfrm_wdat[0]) );
  INVX1 U139 ( .A(n44), .Y(n191) );
  INVX1 U140 ( .A(hit_xd), .Y(n158) );
  NAND21XL U141 ( .B(esfrm_oe), .A(n219), .Y(esfrm_rrdy) );
  MUX2X1 U142 ( .D0(n180), .D1(n176), .S(bist_en), .Y(iram_ce) );
  OAI211X1 U143 ( .C(n165), .D(n176), .A(n3), .B(n175), .Y(xram_we) );
  OAI222XL U144 ( .A(n167), .B(n166), .C(bist_xram), .D(n165), .E(n164), .F(
        n163), .Y(iram_we) );
  AND2X1 U145 ( .A(n24), .B(n68), .Y(N44) );
  OAI21BBXL U146 ( .A(n40), .B(n39), .C(n156), .Y(n43) );
  INVX1 U147 ( .A(n42), .Y(n171) );
  NAND21XL U148 ( .B(n41), .A(n7), .Y(n42) );
  NAND21X1 U149 ( .B(n10), .A(bist_wdat[6]), .Y(n82) );
  INVX1 U150 ( .A(n160), .Y(n40) );
  INVX1 U151 ( .A(iram_a[9]), .Y(n120) );
  NAND43X1 U152 ( .B(n180), .C(n162), .D(n179), .A(dma_hit_x), .Y(n175) );
  INVX1 U153 ( .A(n202), .Y(n107) );
  OAI32X1 U154 ( .A(n181), .B(n180), .C(n179), .D(xram_rdsel[0]), .E(n178), 
        .Y(dma_ack) );
  INVX1 U155 ( .A(n200), .Y(n150) );
  MUX2XL U156 ( .D0(addr1[1]), .D1(addr0[1]), .S(n104), .Y(esfrm_adr[1]) );
  MUX2XL U157 ( .D0(addr1[2]), .D1(addr0[2]), .S(n104), .Y(esfrm_adr[2]) );
  OAI211X1 U158 ( .C(n90), .D(n126), .A(n132), .B(n89), .Y(xram_a[0]) );
  NOR2X2 U159 ( .A(n17), .B(cpurst), .Y(memack) );
  AOI21X1 U160 ( .B(xram_rdsel[0]), .C(xram_rdsel[1]), .A(n177), .Y(n17) );
  INVXL U161 ( .A(n140), .Y(esfrm_adr[3]) );
  GEN3XL U162 ( .F(xram_rdsel[0]), .G(n178), .E(n154), .D(n31), .C(n181), .B(
        n28), .A(n180), .Y(n44) );
  NAND32X1 U163 ( .B(dma_w), .C(n26), .A(xram_rdsel[0]), .Y(n28) );
  AO21X1 U164 ( .B(n154), .C(n25), .A(xram_rdsel[1]), .Y(n26) );
  INVX1 U165 ( .A(memrd_c), .Y(n25) );
  NAND21X1 U166 ( .B(dma_w), .A(memrd_c), .Y(n31) );
  INVX1 U167 ( .A(n38), .Y(n190) );
  GEN2XL U168 ( .D(xram_rdsel[0]), .E(n37), .C(n41), .B(n36), .A(n35), .Y(n38)
         );
  NAND21X1 U169 ( .B(dma_r), .A(n32), .Y(n36) );
  GEN2XL U170 ( .D(n34), .E(n33), .C(xram_rdsel[1]), .B(n37), .A(n180), .Y(n35) );
  OAI221X1 U171 ( .A(n167), .B(n148), .C(n164), .D(n151), .E(n147), .Y(
        iram_a[7]) );
  OAI211X1 U172 ( .C(n148), .D(n126), .A(n147), .B(n113), .Y(xram_a[7]) );
  INVX1 U173 ( .A(r_pg0_sel[0]), .Y(n148) );
  OAI211X1 U174 ( .C(n50), .D(n66), .A(n70), .B(n49), .Y(xram_d[0]) );
  AOI22X1 U175 ( .A(memdatao[0]), .B(n64), .C(dma_wdat[0]), .D(n63), .Y(n49)
         );
  OAI211X1 U176 ( .C(n128), .D(n124), .A(n123), .B(n122), .Y(xram_a[9]) );
  INVX1 U177 ( .A(memaddr[9]), .Y(n124) );
  OA21X1 U178 ( .B(n131), .C(n121), .A(n120), .Y(n122) );
  NAND21X1 U179 ( .B(n45), .A(xram_rdsel[1]), .Y(n37) );
  AOI222XL U180 ( .A(dma_addr[7]), .B(n112), .C(n111), .D(n110), .E(n118), .F(
        n109), .Y(n113) );
  OAI31XL U181 ( .A(n200), .B(memaddr[10]), .C(n107), .D(n106), .Y(n110) );
  OAI31XL U182 ( .A(n200), .B(n108), .C(memaddr_c[10]), .D(n199), .Y(n109) );
  OA222X1 U183 ( .A(n128), .B(n201), .C(n127), .D(n126), .E(n194), .F(n125), 
        .Y(n129) );
  OA222X1 U184 ( .A(n131), .B(n116), .C(n115), .D(n125), .E(n128), .F(n114), 
        .Y(n117) );
  INVX1 U185 ( .A(dma_addr[8]), .Y(n116) );
  INVX1 U186 ( .A(memaddr[8]), .Y(n114) );
  INVX1 U187 ( .A(memaddr_c[8]), .Y(n115) );
  AOI32X1 U188 ( .A(n119), .B(r_pg0_sel[2]), .C(n187), .D(n118), .E(
        memaddr_c[9]), .Y(n123) );
  INVX1 U189 ( .A(esfrm_wdat[1]), .Y(n52) );
  AOI22X1 U190 ( .A(memdatao[1]), .B(n64), .C(dma_wdat[1]), .D(n63), .Y(n51)
         );
  AO21X1 U191 ( .B(r_pg0_sel[1]), .C(n19), .A(n6), .Y(n160) );
  NAND2X1 U192 ( .A(n187), .B(r_pg0_sel[3]), .Y(n127) );
  OAI211X1 U193 ( .C(r_pg0_sel[1]), .D(r_pg0_sel[0]), .A(r_pg0_sel[2]), .B(
        r_pg0_sel[3]), .Y(n187) );
  OAI211X1 U194 ( .C(n58), .D(n66), .A(n78), .B(n57), .Y(xram_d[4]) );
  INVX1 U195 ( .A(esfrm_wdat[4]), .Y(n58) );
  AOI22X1 U196 ( .A(memdatao[4]), .B(n64), .C(dma_wdat[4]), .D(n63), .Y(n57)
         );
  OAI211X1 U197 ( .C(n60), .D(n66), .A(n80), .B(n59), .Y(xram_d[5]) );
  INVX1 U198 ( .A(esfrm_wdat[5]), .Y(n60) );
  AOI22X1 U199 ( .A(memdatao[5]), .B(n64), .C(dma_wdat[5]), .D(n63), .Y(n59)
         );
  OAI211X1 U200 ( .C(n54), .D(n66), .A(n74), .B(n53), .Y(xram_d[2]) );
  INVX1 U201 ( .A(esfrm_wdat[2]), .Y(n54) );
  AOI22X1 U202 ( .A(memdatao[2]), .B(n64), .C(dma_wdat[2]), .D(n63), .Y(n53)
         );
  OAI211X1 U203 ( .C(n56), .D(n66), .A(n76), .B(n55), .Y(xram_d[3]) );
  INVX1 U204 ( .A(esfrm_wdat[3]), .Y(n56) );
  AOI22X1 U205 ( .A(memdatao[3]), .B(n64), .C(dma_wdat[3]), .D(n63), .Y(n55)
         );
  OAI211X1 U206 ( .C(n67), .D(n66), .A(n84), .B(n65), .Y(xram_d[7]) );
  INVX1 U207 ( .A(esfrm_wdat[7]), .Y(n67) );
  AOI22X1 U208 ( .A(memdatao[7]), .B(n64), .C(dma_wdat[7]), .D(n63), .Y(n65)
         );
  OAI211X1 U209 ( .C(n62), .D(n66), .A(n82), .B(n61), .Y(xram_d[6]) );
  INVX1 U210 ( .A(esfrm_wdat[6]), .Y(n62) );
  AOI22X1 U211 ( .A(memdatao[6]), .B(n64), .C(dma_wdat[6]), .D(n63), .Y(n61)
         );
  INVX1 U212 ( .A(r_i2c_attr), .Y(n186) );
  AO222X1 U213 ( .A(xram_rdat[7]), .B(n40), .C(iram_rdat[7]), .D(n30), .E(
        regx_rdat[7]), .F(n7), .Y(n221) );
  NOR2X1 U214 ( .A(delay_rrdy), .B(r_pg0_rdrdy), .Y(n219) );
  AO222X1 U215 ( .A(xram_rdat[1]), .B(n40), .C(iram_rdat[1]), .D(n30), .E(
        regx_rdat[1]), .F(n7), .Y(n227) );
  AO222X1 U216 ( .A(xram_rdat[4]), .B(n40), .C(iram_rdat[4]), .D(n30), .E(
        regx_rdat[4]), .F(n7), .Y(n224) );
  INVX1 U217 ( .A(idat_adr[7]), .Y(n151) );
  AO222X1 U218 ( .A(xram_rdat[2]), .B(n40), .C(iram_rdat[2]), .D(n30), .E(
        regx_rdat[2]), .F(n7), .Y(n226) );
  AO222X1 U219 ( .A(xram_rdat[3]), .B(n40), .C(iram_rdat[3]), .D(n30), .E(
        regx_rdat[3]), .F(n7), .Y(n225) );
  AO222X1 U220 ( .A(xram_rdat[5]), .B(n40), .C(iram_rdat[5]), .D(n30), .E(
        regx_rdat[5]), .F(n7), .Y(n223) );
  AO222X1 U221 ( .A(xram_rdat[6]), .B(n40), .C(iram_rdat[6]), .D(n8), .E(
        regx_rdat[6]), .F(n7), .Y(n222) );
  AO222X1 U222 ( .A(xram_rdat[0]), .B(n40), .C(iram_rdat[0]), .D(n8), .E(
        regx_rdat[0]), .F(n7), .Y(n228) );
  INVX1 U223 ( .A(xram_rdsel[0]), .Y(n33) );
  NAND21X1 U224 ( .B(n9), .A(bist_adr[3]), .Y(n139) );
  NAND21X1 U225 ( .B(n9), .A(bist_adr[5]), .Y(n143) );
  NAND21X1 U226 ( .B(n9), .A(bist_adr[2]), .Y(n137) );
  NAND21X1 U227 ( .B(n9), .A(bist_adr[1]), .Y(n134) );
  NAND21X1 U228 ( .B(n9), .A(bist_adr[0]), .Y(n132) );
  NAND21X1 U229 ( .B(n9), .A(bist_adr[6]), .Y(n144) );
  NAND21X1 U230 ( .B(n9), .A(bist_adr[4]), .Y(n141) );
  OR2X1 U231 ( .A(memrd), .B(memwr), .Y(n87) );
  NAND21X1 U232 ( .B(n9), .A(bist_wdat[7]), .Y(n84) );
  NAND21X1 U233 ( .B(n10), .A(bist_adr[7]), .Y(n147) );
  NAND21X1 U234 ( .B(n10), .A(bist_adr[10]), .Y(n152) );
  INVX1 U235 ( .A(memaddr[7]), .Y(n106) );
  INVX1 U236 ( .A(xram_rdsel[1]), .Y(n178) );
  INVX1 U237 ( .A(dma_w), .Y(n179) );
  INVX1 U238 ( .A(dma_r), .Y(n154) );
  INVX1 U239 ( .A(bist_xram), .Y(n176) );
  INVX1 U240 ( .A(dma_addr[10]), .Y(n130) );
  INVX1 U241 ( .A(dma_addr[9]), .Y(n121) );
  MUX2IX2 U242 ( .D0(addr1[7]), .D1(addr0[7]), .S(n104), .Y(n183) );
  MUX2XL U243 ( .D0(wdat0[2]), .D1(wdat1[2]), .S(i_wr[1]), .Y(esfrm_wdat[2])
         );
  MUX2XL U244 ( .D0(wdat0[7]), .D1(wdat1[7]), .S(i_wr[1]), .Y(esfrm_wdat[7])
         );
  MUX2XL U245 ( .D0(wdat0[1]), .D1(wdat1[1]), .S(i_wr[1]), .Y(esfrm_wdat[1])
         );
  MUX2XL U246 ( .D0(wdat0[3]), .D1(wdat1[3]), .S(i_wr[1]), .Y(esfrm_wdat[3])
         );
  NAND21XL U247 ( .B(n30), .A(n29), .Y(n47) );
  AO21XL U248 ( .B(n40), .C(n29), .A(n27), .Y(n24) );
  AND2XL U249 ( .A(n189), .B(n188), .Y(sfrack) );
  INVX2 U250 ( .A(n183), .Y(n184) );
  NAND32X1 U251 ( .B(n27), .C(n68), .A(n156), .Y(n180) );
  INVX2 U252 ( .A(n189), .Y(esfrm_we) );
  OAI211X1 U253 ( .C(n187), .D(n186), .A(n185), .B(n184), .Y(n189) );
  MUX2IXL U254 ( .D0(wdat0[0]), .D1(wdat1[0]), .S(i_wr[1]), .Y(n50) );
  MUX2XL U255 ( .D0(wdat0[5]), .D1(wdat1[5]), .S(i_wr[1]), .Y(esfrm_wdat[5])
         );
  MUX2XL U256 ( .D0(wdat0[6]), .D1(wdat1[6]), .S(i_wr[1]), .Y(esfrm_wdat[6])
         );
  MUX2XL U257 ( .D0(wdat0[4]), .D1(wdat1[4]), .S(i_wr[1]), .Y(esfrm_wdat[4])
         );
  AO222XL U258 ( .A(delay_rdat[7]), .B(n220), .C(r_pg0_rdrdy), .D(n221), .E(
        mcu_esfr_rdat[7]), .F(n219), .Y(esfrm_rdat[7]) );
  NAND21XL U259 ( .B(n192), .A(n155), .Y(n162) );
  NAND6X2 U260 ( .A(memwr), .B(n166), .C(n156), .D(n155), .E(n154), .F(n179), 
        .Y(n159) );
  AOI222XL U261 ( .A(memaddr[6]), .B(n111), .C(n119), .D(esfrm_adr[6]), .E(
        memaddr_c[6]), .F(n118), .Y(n105) );
  AOI222XL U262 ( .A(dma_addr[0]), .B(n112), .C(memaddr_c[0]), .D(n118), .E(
        memaddr[0]), .F(n111), .Y(n89) );
  AOI222XL U263 ( .A(memaddr[1]), .B(n111), .C(n119), .D(esfrm_adr[1]), .E(
        memaddr_c[1]), .F(n118), .Y(n91) );
  AO222XL U264 ( .A(delay_rdat[1]), .B(n220), .C(r_pg0_rdrdy), .D(n227), .E(
        mcu_esfr_rdat[1]), .F(n219), .Y(esfrm_rdat[1]) );
  AOI222XL U265 ( .A(memaddr[4]), .B(n111), .C(n119), .D(esfrm_adr[4]), .E(
        memaddr_c[4]), .F(n118), .Y(n98) );
  MUX2IXL U266 ( .D0(addr1[4]), .D1(addr0[4]), .S(n104), .Y(n142) );
  MUX2IXL U267 ( .D0(addr1[3]), .D1(addr0[3]), .S(n104), .Y(n140) );
  MUX2IXL U268 ( .D0(addr1[0]), .D1(addr0[0]), .S(n104), .Y(n90) );
  MUX2IXL U269 ( .D0(addr1[6]), .D1(addr0[6]), .S(n104), .Y(n146) );
  AO222XL U270 ( .A(delay_rdat[4]), .B(n220), .C(r_pg0_rdrdy), .D(n224), .E(
        mcu_esfr_rdat[4]), .F(n219), .Y(esfrm_rdat[4]) );
  AOI222XL U271 ( .A(memaddr[2]), .B(n111), .C(n119), .D(esfrm_adr[2]), .E(
        memaddr_c[2]), .F(n118), .Y(n92) );
  OAI21X1 U272 ( .B(dma_addr[9]), .C(dma_addr[8]), .A(dma_addr[10]), .Y(
        dma_hit_x) );
  OAI21X1 U273 ( .B(n194), .C(n195), .A(n196), .Y(n193) );
  INVX1 U274 ( .A(r_pg0_sel[1]), .Y(n197) );
  NAND4X1 U275 ( .A(memaddr_c[14]), .B(memaddr_c[13]), .C(memaddr_c[15]), .D(
        n204), .Y(n203) );
  NOR32XL U276 ( .B(memaddr_c[12]), .C(memaddr_c[11]), .A(n199), .Y(n204) );
  NOR21XL U277 ( .B(bist_adr[9]), .A(n10), .Y(iram_a[9]) );
  INVX1 U278 ( .A(bist_adr[8]), .Y(n198) );
  INVX1 U279 ( .A(channel_sel), .Y(n200) );
  MUX2IX1 U280 ( .D0(n209), .D1(n210), .S(idat_adr[6]), .Y(n208) );
  NAND2X1 U281 ( .A(idat_adr[4]), .B(idat_adr[5]), .Y(n210) );
  AOI21X1 U282 ( .B(n207), .C(n206), .A(n205), .Y(n209) );
  INVX1 U283 ( .A(idat_adr[5]), .Y(n205) );
  INVX1 U284 ( .A(idat_adr[4]), .Y(n206) );
  INVX1 U285 ( .A(idat_adr[3]), .Y(n207) );
  NOR43XL U286 ( .B(memaddr[15]), .C(memaddr[13]), .D(memaddr[14]), .A(n213), 
        .Y(n212) );
  NOR32XL U287 ( .B(memaddr[8]), .C(memaddr[9]), .A(n201), .Y(n211) );
  NOR4XL U288 ( .A(memaddr[14]), .B(memaddr[15]), .C(memaddr[13]), .D(n214), 
        .Y(hit_xd) );
  OAI211X1 U289 ( .C(n201), .D(n202), .A(n213), .B(n215), .Y(n214) );
  INVX1 U290 ( .A(memaddr[12]), .Y(n213) );
  AOI211X1 U291 ( .C(memaddr_c[14]), .D(n216), .A(memaddr_c[15]), .B(cpurst), 
        .Y(hit_ps_c) );
  NAND4X1 U292 ( .A(n195), .B(n196), .C(n194), .D(n199), .Y(n216) );
  INVX1 U293 ( .A(memaddr_c[7]), .Y(n199) );
  INVX1 U294 ( .A(memaddr_c[10]), .Y(n194) );
  NOR3XL U295 ( .A(memaddr_c[12]), .B(memaddr_c[13]), .C(memaddr_c[11]), .Y(
        n196) );
  NOR2X1 U296 ( .A(memaddr_c[8]), .B(memaddr_c[9]), .Y(n195) );
  AOI211X1 U297 ( .C(memaddr[14]), .D(n217), .A(memaddr[15]), .B(cpurst), .Y(
        hit_ps) );
  NAND4X1 U298 ( .A(n201), .B(n215), .C(n202), .D(n218), .Y(n217) );
  NOR3XL U299 ( .A(memaddr[12]), .B(memaddr[7]), .C(memaddr[13]), .Y(n218) );
  NOR2X1 U300 ( .A(memaddr[8]), .B(memaddr[9]), .Y(n202) );
  INVX1 U301 ( .A(memaddr[11]), .Y(n215) );
  INVX1 U302 ( .A(memaddr[10]), .Y(n201) );
  AO222X1 U303 ( .A(delay_rdat[6]), .B(n220), .C(r_pg0_rdrdy), .D(n222), .E(
        mcu_esfr_rdat[6]), .F(n219), .Y(esfrm_rdat[6]) );
  AO222X1 U304 ( .A(delay_rdat[5]), .B(n220), .C(r_pg0_rdrdy), .D(n223), .E(
        mcu_esfr_rdat[5]), .F(n219), .Y(esfrm_rdat[5]) );
  AO222X1 U305 ( .A(delay_rdat[3]), .B(n220), .C(r_pg0_rdrdy), .D(n225), .E(
        mcu_esfr_rdat[3]), .F(n219), .Y(esfrm_rdat[3]) );
  AO222X1 U306 ( .A(delay_rdat[2]), .B(n220), .C(r_pg0_rdrdy), .D(n226), .E(
        mcu_esfr_rdat[2]), .F(n219), .Y(esfrm_rdat[2]) );
  AO222X1 U307 ( .A(delay_rdat[0]), .B(n220), .C(r_pg0_rdrdy), .D(n228), .E(
        mcu_esfr_rdat[0]), .F(n219), .Y(esfrm_rdat[0]) );
  NOR21XL U308 ( .B(delay_rrdy), .A(r_pg0_rdrdy), .Y(n220) );
endmodule

